`include "parameter.v"

(*DONT_TOUCH = "true"*)
module tf_ROM (
input clk,
input [`ADDR_ROM_WIDTH-1:0] A,
input REN,
output reg [`P*`DATA_WIDTH-1:0] Q //同时给出 P 个 twiddle factor
);
/*
基4修改：同时输出多个twiddle向量。
radix-4：Q = {W1_vec, W2_vec, W3_vec}（多组打包）
*/

// (*rom_style = "block"*) reg [`P*`DATA_WIDTH-1:0] bank [`ROM_DEPTH-1:0];

// always@(posedge clk)
// begin
//     if(REN == 1'b1) 
//         Q <= bank[A];
//     else
//         Q <='b0;
// end

`ifdef OP0
    always@(posedge clk)
        begin
        if(REN == 1'b1) begin
        case(A)
        10'd0:   Q <= 24'b011011000001011011000001;
        10'd1:   Q <= 24'b011011000001011011000001;
        10'd2:   Q <= 24'b011011000001011011000001;
        10'd3:   Q <= 24'b011011000001011011000001;
        10'd4:   Q <= 24'b011011000001011011000001;
        10'd5:   Q <= 24'b011011000001011011000001;
        10'd6:   Q <= 24'b011011000001011011000001;
        10'd7:   Q <= 24'b011011000001011011000001;
        10'd8:   Q <= 24'b011011000001011011000001;
        10'd9:   Q <= 24'b011011000001011011000001;
        10'd10:  Q <= 24'b011011000001011011000001;
        10'd11:  Q <= 24'b011011000001011011000001;
        10'd12:  Q <= 24'b011011000001011011000001;
        10'd13:  Q <= 24'b011011000001011011000001;
        10'd14:  Q <= 24'b011011000001011011000001;
        10'd15:  Q <= 24'b011011000001011011000001;
        10'd16:  Q <= 24'b011011000001011011000001;
        10'd17:  Q <= 24'b011011000001011011000001;
        10'd18:  Q <= 24'b011011000001011011000001;
        10'd19:  Q <= 24'b011011000001011011000001;
        10'd20:  Q <= 24'b011011000001011011000001;
        10'd21:  Q <= 24'b011011000001011011000001;
        10'd22:  Q <= 24'b011011000001011011000001;
        10'd23:  Q <= 24'b011011000001011011000001;
        10'd24:  Q <= 24'b011011000001011011000001;
        10'd25:  Q <= 24'b011011000001011011000001;
        10'd26:  Q <= 24'b011011000001011011000001;
        10'd27:  Q <= 24'b011011000001011011000001;
        10'd28:  Q <= 24'b011011000001011011000001;
        10'd29:  Q <= 24'b011011000001011011000001;
        10'd30:  Q <= 24'b011011000001011011000001;
        10'd31:  Q <= 24'b011011000001011011000001;
        10'd32:  Q <= 24'b011011000001011011000001;
        10'd33:  Q <= 24'b011011000001011011000001;
        10'd34:  Q <= 24'b011011000001011011000001;
        10'd35:  Q <= 24'b011011000001011011000001;
        10'd36:  Q <= 24'b011011000001011011000001;
        10'd37:  Q <= 24'b011011000001011011000001;
        10'd38:  Q <= 24'b011011000001011011000001;
        10'd39:  Q <= 24'b011011000001011011000001;
        10'd40:  Q <= 24'b011011000001011011000001;
        10'd41:  Q <= 24'b011011000001011011000001;
        10'd42:  Q <= 24'b011011000001011011000001;
        10'd43:  Q <= 24'b011011000001011011000001;
        10'd44:  Q <= 24'b011011000001011011000001;
        10'd45:  Q <= 24'b011011000001011011000001;
        10'd46:  Q <= 24'b011011000001011011000001;
        10'd47:  Q <= 24'b011011000001011011000001;
        10'd48:  Q <= 24'b011011000001011011000001;
        10'd49:  Q <= 24'b011011000001011011000001;
        10'd50:  Q <= 24'b011011000001011011000001;
        10'd51:  Q <= 24'b011011000001011011000001;
        10'd52:  Q <= 24'b011011000001011011000001;
        10'd53:  Q <= 24'b011011000001011011000001;
        10'd54:  Q <= 24'b011011000001011011000001;
        10'd55:  Q <= 24'b011011000001011011000001;
        10'd56:  Q <= 24'b011011000001011011000001;
        10'd57:  Q <= 24'b011011000001011011000001;
        10'd58:  Q <= 24'b011011000001011011000001;
        10'd59:  Q <= 24'b011011000001011011000001;
        10'd60:  Q <= 24'b011011000001011011000001;
        10'd61:  Q <= 24'b011011000001011011000001;
        10'd62:  Q <= 24'b011011000001011011000001;
        10'd63:  Q <= 24'b011011000001011011000001;
        10'd64:  Q <= 24'b101000010100101000010100;
        10'd65:  Q <= 24'b101000010100101000010100;
        10'd66:  Q <= 24'b101000010100101000010100;
        10'd67:  Q <= 24'b101000010100101000010100;
        10'd68:  Q <= 24'b101000010100101000010100;
        10'd69:  Q <= 24'b101000010100101000010100;
        10'd70:  Q <= 24'b101000010100101000010100;
        10'd71:  Q <= 24'b101000010100101000010100;
        10'd72:  Q <= 24'b101000010100101000010100;
        10'd73:  Q <= 24'b101000010100101000010100;
        10'd74:  Q <= 24'b101000010100101000010100;
        10'd75:  Q <= 24'b101000010100101000010100;
        10'd76:  Q <= 24'b101000010100101000010100;
        10'd77:  Q <= 24'b101000010100101000010100;
        10'd78:  Q <= 24'b101000010100101000010100;
        10'd79:  Q <= 24'b101000010100101000010100;
        10'd80:  Q <= 24'b101000010100101000010100;
        10'd81:  Q <= 24'b101000010100101000010100;
        10'd82:  Q <= 24'b101000010100101000010100;
        10'd83:  Q <= 24'b101000010100101000010100;
        10'd84:  Q <= 24'b101000010100101000010100;
        10'd85:  Q <= 24'b101000010100101000010100;
        10'd86:  Q <= 24'b101000010100101000010100;
        10'd87:  Q <= 24'b101000010100101000010100;
        10'd88:  Q <= 24'b101000010100101000010100;
        10'd89:  Q <= 24'b101000010100101000010100;
        10'd90:  Q <= 24'b101000010100101000010100;
        10'd91:  Q <= 24'b101000010100101000010100;
        10'd92:  Q <= 24'b101000010100101000010100;
        10'd93:  Q <= 24'b101000010100101000010100;
        10'd94:  Q <= 24'b101000010100101000010100;
        10'd95:  Q <= 24'b101000010100101000010100;
        10'd96:  Q <= 24'b110011011001110011011001;
        10'd97:  Q <= 24'b110011011001110011011001;
        10'd98:  Q <= 24'b110011011001110011011001;
        10'd99:  Q <= 24'b110011011001110011011001;
        10'd100: Q <= 24'b110011011001110011011001;
        10'd101: Q <= 24'b110011011001110011011001;
        10'd102: Q <= 24'b110011011001110011011001;
        10'd103: Q <= 24'b110011011001110011011001;
        10'd104: Q <= 24'b110011011001110011011001;
        10'd105: Q <= 24'b110011011001110011011001;
        10'd106: Q <= 24'b110011011001110011011001;
        10'd107: Q <= 24'b110011011001110011011001;
        10'd108: Q <= 24'b110011011001110011011001;
        10'd109: Q <= 24'b110011011001110011011001;
        10'd110: Q <= 24'b110011011001110011011001;
        10'd111: Q <= 24'b110011011001110011011001;
        10'd112: Q <= 24'b110011011001110011011001;
        10'd113: Q <= 24'b110011011001110011011001;
        10'd114: Q <= 24'b110011011001110011011001;
        10'd115: Q <= 24'b110011011001110011011001;
        10'd116: Q <= 24'b110011011001110011011001;
        10'd117: Q <= 24'b110011011001110011011001;
        10'd118: Q <= 24'b110011011001110011011001;
        10'd119: Q <= 24'b110011011001110011011001;
        10'd120: Q <= 24'b110011011001110011011001;
        10'd121: Q <= 24'b110011011001110011011001;
        10'd122: Q <= 24'b110011011001110011011001;
        10'd123: Q <= 24'b110011011001110011011001;
        10'd124: Q <= 24'b110011011001110011011001;
        10'd125: Q <= 24'b110011011001110011011001;
        10'd126: Q <= 24'b110011011001110011011001;
        10'd127: Q <= 24'b110011011001110011011001;
        10'd128: Q <= 24'b101001010010101001010010;
        10'd129: Q <= 24'b101001010010101001010010;
        10'd130: Q <= 24'b101001010010101001010010;
        10'd131: Q <= 24'b101001010010101001010010;
        10'd132: Q <= 24'b101001010010101001010010;
        10'd133: Q <= 24'b101001010010101001010010;
        10'd134: Q <= 24'b101001010010101001010010;
        10'd135: Q <= 24'b101001010010101001010010;
        10'd136: Q <= 24'b101001010010101001010010;
        10'd137: Q <= 24'b101001010010101001010010;
        10'd138: Q <= 24'b101001010010101001010010;
        10'd139: Q <= 24'b101001010010101001010010;
        10'd140: Q <= 24'b101001010010101001010010;
        10'd141: Q <= 24'b101001010010101001010010;
        10'd142: Q <= 24'b101001010010101001010010;
        10'd143: Q <= 24'b101001010010101001010010;
        10'd144: Q <= 24'b001001110110001001110110;
        10'd145: Q <= 24'b001001110110001001110110;
        10'd146: Q <= 24'b001001110110001001110110;
        10'd147: Q <= 24'b001001110110001001110110;
        10'd148: Q <= 24'b001001110110001001110110;
        10'd149: Q <= 24'b001001110110001001110110;
        10'd150: Q <= 24'b001001110110001001110110;
        10'd151: Q <= 24'b001001110110001001110110;
        10'd152: Q <= 24'b001001110110001001110110;
        10'd153: Q <= 24'b001001110110001001110110;
        10'd154: Q <= 24'b001001110110001001110110;
        10'd155: Q <= 24'b001001110110001001110110;
        10'd156: Q <= 24'b001001110110001001110110;
        10'd157: Q <= 24'b001001110110001001110110;
        10'd158: Q <= 24'b001001110110001001110110;
        10'd159: Q <= 24'b001001110110001001110110;
        10'd160: Q <= 24'b011101101001011101101001;
        10'd161: Q <= 24'b011101101001011101101001;
        10'd162: Q <= 24'b011101101001011101101001;
        10'd163: Q <= 24'b011101101001011101101001;
        10'd164: Q <= 24'b011101101001011101101001;
        10'd165: Q <= 24'b011101101001011101101001;
        10'd166: Q <= 24'b011101101001011101101001;
        10'd167: Q <= 24'b011101101001011101101001;
        10'd168: Q <= 24'b011101101001011101101001;
        10'd169: Q <= 24'b011101101001011101101001;
        10'd170: Q <= 24'b011101101001011101101001;
        10'd171: Q <= 24'b011101101001011101101001;
        10'd172: Q <= 24'b011101101001011101101001;
        10'd173: Q <= 24'b011101101001011101101001;
        10'd174: Q <= 24'b011101101001011101101001;
        10'd175: Q <= 24'b011101101001011101101001;
        10'd176: Q <= 24'b001101010000001101010000;
        10'd177: Q <= 24'b001101010000001101010000;
        10'd178: Q <= 24'b001101010000001101010000;
        10'd179: Q <= 24'b001101010000001101010000;
        10'd180: Q <= 24'b001101010000001101010000;
        10'd181: Q <= 24'b001101010000001101010000;
        10'd182: Q <= 24'b001101010000001101010000;
        10'd183: Q <= 24'b001101010000001101010000;
        10'd184: Q <= 24'b001101010000001101010000;
        10'd185: Q <= 24'b001101010000001101010000;
        10'd186: Q <= 24'b001101010000001101010000;
        10'd187: Q <= 24'b001101010000001101010000;
        10'd188: Q <= 24'b001101010000001101010000;
        10'd189: Q <= 24'b001101010000001101010000;
        10'd190: Q <= 24'b001101010000001101010000;
        10'd191: Q <= 24'b001101010000001101010000;
        10'd192: Q <= 24'b010000100110010000100110;
        10'd193: Q <= 24'b010000100110010000100110;
        10'd194: Q <= 24'b010000100110010000100110;
        10'd195: Q <= 24'b010000100110010000100110;
        10'd196: Q <= 24'b010000100110010000100110;
        10'd197: Q <= 24'b010000100110010000100110;
        10'd198: Q <= 24'b010000100110010000100110;
        10'd199: Q <= 24'b010000100110010000100110;
        10'd200: Q <= 24'b011101111111011101111111;
        10'd201: Q <= 24'b011101111111011101111111;
        10'd202: Q <= 24'b011101111111011101111111;
        10'd203: Q <= 24'b011101111111011101111111;
        10'd204: Q <= 24'b011101111111011101111111;
        10'd205: Q <= 24'b011101111111011101111111;
        10'd206: Q <= 24'b011101111111011101111111;
        10'd207: Q <= 24'b011101111111011101111111;
        10'd208: Q <= 24'b000011000001000011000001;
        10'd209: Q <= 24'b000011000001000011000001;
        10'd210: Q <= 24'b000011000001000011000001;
        10'd211: Q <= 24'b000011000001000011000001;
        10'd212: Q <= 24'b000011000001000011000001;
        10'd213: Q <= 24'b000011000001000011000001;
        10'd214: Q <= 24'b000011000001000011000001;
        10'd215: Q <= 24'b000011000001000011000001;
        10'd216: Q <= 24'b001100011101001100011101;
        10'd217: Q <= 24'b001100011101001100011101;
        10'd218: Q <= 24'b001100011101001100011101;
        10'd219: Q <= 24'b001100011101001100011101;
        10'd220: Q <= 24'b001100011101001100011101;
        10'd221: Q <= 24'b001100011101001100011101;
        10'd222: Q <= 24'b001100011101001100011101;
        10'd223: Q <= 24'b001100011101001100011101;
        10'd224: Q <= 24'b101011100010101011100010;
        10'd225: Q <= 24'b101011100010101011100010;
        10'd226: Q <= 24'b101011100010101011100010;
        10'd227: Q <= 24'b101011100010101011100010;
        10'd228: Q <= 24'b101011100010101011100010;
        10'd229: Q <= 24'b101011100010101011100010;
        10'd230: Q <= 24'b101011100010101011100010;
        10'd231: Q <= 24'b101011100010101011100010;
        10'd232: Q <= 24'b110010111100110010111100;
        10'd233: Q <= 24'b110010111100110010111100;
        10'd234: Q <= 24'b110010111100110010111100;
        10'd235: Q <= 24'b110010111100110010111100;
        10'd236: Q <= 24'b110010111100110010111100;
        10'd237: Q <= 24'b110010111100110010111100;
        10'd238: Q <= 24'b110010111100110010111100;
        10'd239: Q <= 24'b110010111100110010111100;
        10'd240: Q <= 24'b001000111001001000111001;
        10'd241: Q <= 24'b001000111001001000111001;
        10'd242: Q <= 24'b001000111001001000111001;
        10'd243: Q <= 24'b001000111001001000111001;
        10'd244: Q <= 24'b001000111001001000111001;
        10'd245: Q <= 24'b001000111001001000111001;
        10'd246: Q <= 24'b001000111001001000111001;
        10'd247: Q <= 24'b001000111001001000111001;
        10'd248: Q <= 24'b011011010010011011010010;
        10'd249: Q <= 24'b011011010010011011010010;
        10'd250: Q <= 24'b011011010010011011010010;
        10'd251: Q <= 24'b011011010010011011010010;
        10'd252: Q <= 24'b011011010010011011010010;
        10'd253: Q <= 24'b011011010010011011010010;
        10'd254: Q <= 24'b011011010010011011010010;
        10'd255: Q <= 24'b011011010010011011010010;
        10'd256: Q <= 24'b000100101000000100101000;
        10'd257: Q <= 24'b000100101000000100101000;
        10'd258: Q <= 24'b000100101000000100101000;
        10'd259: Q <= 24'b000100101000000100101000;
        10'd260: Q <= 24'b100110001111100110001111;
        10'd261: Q <= 24'b100110001111100110001111;
        10'd262: Q <= 24'b100110001111100110001111;
        10'd263: Q <= 24'b100110001111100110001111;
        10'd264: Q <= 24'b010100111011010100111011;
        10'd265: Q <= 24'b010100111011010100111011;
        10'd266: Q <= 24'b010100111011010100111011;
        10'd267: Q <= 24'b010100111011010100111011;
        10'd268: Q <= 24'b010111000100010111000100;
        10'd269: Q <= 24'b010111000100010111000100;
        10'd270: Q <= 24'b010111000100010111000100;
        10'd271: Q <= 24'b010111000100010111000100;
        10'd272: Q <= 24'b101111100110101111100110;
        10'd273: Q <= 24'b101111100110101111100110;
        10'd274: Q <= 24'b101111100110101111100110;
        10'd275: Q <= 24'b101111100110101111100110;
        10'd276: Q <= 24'b000000111000000000111000;
        10'd277: Q <= 24'b000000111000000000111000;
        10'd278: Q <= 24'b000000111000000000111000;
        10'd279: Q <= 24'b000000111000000000111000;
        10'd280: Q <= 24'b100011000000100011000000;
        10'd281: Q <= 24'b100011000000100011000000;
        10'd282: Q <= 24'b100011000000100011000000;
        10'd283: Q <= 24'b100011000000100011000000;
        10'd284: Q <= 24'b010100110101010100110101;
        10'd285: Q <= 24'b010100110101010100110101;
        10'd286: Q <= 24'b010100110101010100110101;
        10'd287: Q <= 24'b010100110101010100110101;
        10'd288: Q <= 24'b010110010010010110010010;
        10'd289: Q <= 24'b010110010010010110010010;
        10'd290: Q <= 24'b010110010010010110010010;
        10'd291: Q <= 24'b010110010010010110010010;
        10'd292: Q <= 24'b100000101110100000101110;
        10'd293: Q <= 24'b100000101110100000101110;
        10'd294: Q <= 24'b100000101110100000101110;
        10'd295: Q <= 24'b100000101110100000101110;
        10'd296: Q <= 24'b001000010111001000010111;
        10'd297: Q <= 24'b001000010111001000010111;
        10'd298: Q <= 24'b001000010111001000010111;
        10'd299: Q <= 24'b001000010111001000010111;
        10'd300: Q <= 24'b101101000010101101000010;
        10'd301: Q <= 24'b101101000010101101000010;
        10'd302: Q <= 24'b101101000010101101000010;
        10'd303: Q <= 24'b101101000010101101000010;
        10'd304: Q <= 24'b100101011001100101011001;
        10'd305: Q <= 24'b100101011001100101011001;
        10'd306: Q <= 24'b100101011001100101011001;
        10'd307: Q <= 24'b100101011001100101011001;
        10'd308: Q <= 24'b101100111111101100111111;
        10'd309: Q <= 24'b101100111111101100111111;
        10'd310: Q <= 24'b101100111111101100111111;
        10'd311: Q <= 24'b101100111111101100111111;
        10'd312: Q <= 24'b011110110110011110110110;
        10'd313: Q <= 24'b011110110110011110110110;
        10'd314: Q <= 24'b011110110110011110110110;
        10'd315: Q <= 24'b011110110110011110110110;
        10'd316: Q <= 24'b001100110101001100110101;
        10'd317: Q <= 24'b001100110101001100110101;
        10'd318: Q <= 24'b001100110101001100110101;
        10'd319: Q <= 24'b001100110101001100110101;
        10'd320: Q <= 24'b000100100001000100100001;
        10'd321: Q <= 24'b000100100001000100100001;
        10'd322: Q <= 24'b000101001011000101001011;
        10'd323: Q <= 24'b000101001011000101001011;
        10'd324: Q <= 24'b110010110101110010110101;
        10'd325: Q <= 24'b110010110101110010110101;
        10'd326: Q <= 24'b011011011100011011011100;
        10'd327: Q <= 24'b011011011100011011011100;
        10'd328: Q <= 24'b010010101101010010101101;
        10'd329: Q <= 24'b010010101101010010101101;
        10'd330: Q <= 24'b100100000000100100000000;
        10'd331: Q <= 24'b100100000000100100000000;
        10'd332: Q <= 24'b100011100101100011100101;
        10'd333: Q <= 24'b100011100101100011100101;
        10'd334: Q <= 24'b100000000111100000000111;
        10'd335: Q <= 24'b100000000111100000000111;
        10'd336: Q <= 24'b001010001010001010001010;
        10'd337: Q <= 24'b001010001010001010001010;
        10'd338: Q <= 24'b011110111001011110111001;
        10'd339: Q <= 24'b011110111001011110111001;
        10'd340: Q <= 24'b100111010001100111010001;
        10'd341: Q <= 24'b100111010001100111010001;
        10'd342: Q <= 24'b001001111000001001111000;
        10'd343: Q <= 24'b001001111000001001111000;
        10'd344: Q <= 24'b101100110001101100110001;
        10'd345: Q <= 24'b101100110001101100110001;
        10'd346: Q <= 24'b000000100001000000100001;
        10'd347: Q <= 24'b000000100001000000100001;
        10'd348: Q <= 24'b010100101000010100101000;
        10'd349: Q <= 24'b010100101000010100101000;
        10'd350: Q <= 24'b011101111011011101111011;
        10'd351: Q <= 24'b011101111011011101111011;
        10'd352: Q <= 24'b100100001111100100001111;
        10'd353: Q <= 24'b100100001111100100001111;
        10'd354: Q <= 24'b010110011011010110011011;
        10'd355: Q <= 24'b010110011011010110011011;
        10'd356: Q <= 24'b001100100111001100100111;
        10'd357: Q <= 24'b001100100111001100100111;
        10'd358: Q <= 24'b000111000100000111000100;
        10'd359: Q <= 24'b000111000100000111000100;
        10'd360: Q <= 24'b010110011110010110011110;
        10'd361: Q <= 24'b010110011110010110011110;
        10'd362: Q <= 24'b101100110100101100110100;
        10'd363: Q <= 24'b101100110100101100110100;
        10'd364: Q <= 24'b010111111110010111111110;
        10'd365: Q <= 24'b010111111110010111111110;
        10'd366: Q <= 24'b100101100010100101100010;
        10'd367: Q <= 24'b100101100010100101100010;
        10'd368: Q <= 24'b101001010111101001010111;
        10'd369: Q <= 24'b101001010111101001010111;
        10'd370: Q <= 24'b101000111001101000111001;
        10'd371: Q <= 24'b101000111001101000111001;
        10'd372: Q <= 24'b010111001001010111001001;
        10'd373: Q <= 24'b010111001001010111001001;
        10'd374: Q <= 24'b001010001000001010001000;
        10'd375: Q <= 24'b001010001000001010001000;
        10'd376: Q <= 24'b100110101010100110101010;
        10'd377: Q <= 24'b100110101010100110101010;
        10'd378: Q <= 24'b110000100110110000100110;
        10'd379: Q <= 24'b110000100110110000100110;
        10'd380: Q <= 24'b010011001011010011001011;
        10'd381: Q <= 24'b010011001011010011001011;
        10'd382: Q <= 24'b001110001110001110001110;
        10'd383: Q <= 24'b001110001110001110001110;
        10'd384: Q <= 24'b000000010001000000010001;
        10'd385: Q <= 24'b101011001001101011001001;
        10'd386: Q <= 24'b001001000111001001000111;
        10'd387: Q <= 24'b101001011001101001011001;
        10'd388: Q <= 24'b011001100101011001100101;
        10'd389: Q <= 24'b001011010011001011010011;
        10'd390: Q <= 24'b100011110000100011110000;
        10'd391: Q <= 24'b010001001100010001001100;
        10'd392: Q <= 24'b010110000001010110000001;
        10'd393: Q <= 24'b101001100110101001100110;
        10'd394: Q <= 24'b110011010001110011010001;
        10'd395: Q <= 24'b000011101001000011101001;
        10'd396: Q <= 24'b001011110100001011110100;
        10'd397: Q <= 24'b100001101100100001101100;
        10'd398: Q <= 24'b101111000111101111000111;
        10'd399: Q <= 24'b101111101010101111101010;
        10'd400: Q <= 24'b011010100111011010100111;
        10'd401: Q <= 24'b011001110011011001110011;
        10'd402: Q <= 24'b101011100101101011100101;
        10'd403: Q <= 24'b011011111101011011111101;
        10'd404: Q <= 24'b011100110111011100110111;
        10'd405: Q <= 24'b001110111000001110111000;
        10'd406: Q <= 24'b010110110101010110110101;
        10'd407: Q <= 24'b101001111111101001111111;
        10'd408: Q <= 24'b001110101011001110101011;
        10'd409: Q <= 24'b100100000100100100000100;
        10'd410: Q <= 24'b100110000101100110000101;
        10'd411: Q <= 24'b100101010100100101010100;
        10'd412: Q <= 24'b001011011101001011011101;
        10'd413: Q <= 24'b100100100001100100100001;
        10'd414: Q <= 24'b000100001100000100001100;
        10'd415: Q <= 24'b001010000001001010000001;
        10'd416: Q <= 24'b011000110000011000110000;
        10'd417: Q <= 24'b100011111010100011111010;
        10'd418: Q <= 24'b011111110101011111110101;
        10'd419: Q <= 24'b110010010100110010010100;
        10'd420: Q <= 24'b000101110111000101110111;
        10'd421: Q <= 24'b100111110101100111110101;
        10'd422: Q <= 24'b100000101010100000101010;
        10'd423: Q <= 24'b011001101101011001101101;
        10'd424: Q <= 24'b010000100111010000100111;
        10'd425: Q <= 24'b000100111111000100111111;
        10'd426: Q <= 24'b101011010101101011010101;
        10'd427: Q <= 24'b001011110101001011110101;
        10'd428: Q <= 24'b100000110011100000110011;
        10'd429: Q <= 24'b001000110001001000110001;
        10'd430: Q <= 24'b100110100010100110100010;
        10'd431: Q <= 24'b101000100010101000100010;
        10'd432: Q <= 24'b101011110100101011110100;
        10'd433: Q <= 24'b010001000100010001000100;
        10'd434: Q <= 24'b000110010011000110010011;
        10'd435: Q <= 24'b010000000010010000000010;
        10'd436: Q <= 24'b010001110111010001110111;
        10'd437: Q <= 24'b100001100110100001100110;
        10'd438: Q <= 24'b101011010111101011010111;
        10'd439: Q <= 24'b001101110110001101110110;
        10'd440: Q <= 24'b011010111010011010111010;
        10'd441: Q <= 24'b010010111100010010111100;
        10'd442: Q <= 24'b011101010010011101010010;
        10'd443: Q <= 24'b010000000101010000000101;
        10'd444: Q <= 24'b100000111110100000111110;
        10'd445: Q <= 24'b101101110111101101110111;
        10'd446: Q <= 24'b001101110101001101110101;
        10'd447: Q <= 24'b100001101010100001101010;
        10'd448: Q <= 24'b011011000001011011000001;
        10'd449: Q <= 24'b011011000001011011000001;
        10'd450: Q <= 24'b011011000001011011000001;
        10'd451: Q <= 24'b011011000001011011000001;
        10'd452: Q <= 24'b011011000001011011000001;
        10'd453: Q <= 24'b011011000001011011000001;
        10'd454: Q <= 24'b011011000001011011000001;
        10'd455: Q <= 24'b011011000001011011000001;
        10'd456: Q <= 24'b011011000001011011000001;
        10'd457: Q <= 24'b011011000001011011000001;
        10'd458: Q <= 24'b011011000001011011000001;
        10'd459: Q <= 24'b011011000001011011000001;
        10'd460: Q <= 24'b011011000001011011000001;
        10'd461: Q <= 24'b011011000001011011000001;
        10'd462: Q <= 24'b011011000001011011000001;
        10'd463: Q <= 24'b011011000001011011000001;
        10'd464: Q <= 24'b011011000001011011000001;
        10'd465: Q <= 24'b011011000001011011000001;
        10'd466: Q <= 24'b011011000001011011000001;
        10'd467: Q <= 24'b011011000001011011000001;
        10'd468: Q <= 24'b011011000001011011000001;
        10'd469: Q <= 24'b011011000001011011000001;
        10'd470: Q <= 24'b011011000001011011000001;
        10'd471: Q <= 24'b011011000001011011000001;
        10'd472: Q <= 24'b011011000001011011000001;
        10'd473: Q <= 24'b011011000001011011000001;
        10'd474: Q <= 24'b011011000001011011000001;
        10'd475: Q <= 24'b011011000001011011000001;
        10'd476: Q <= 24'b011011000001011011000001;
        10'd477: Q <= 24'b011011000001011011000001;
        10'd478: Q <= 24'b011011000001011011000001;
        10'd479: Q <= 24'b011011000001011011000001;
        10'd480: Q <= 24'b011011000001011011000001;
        10'd481: Q <= 24'b011011000001011011000001;
        10'd482: Q <= 24'b011011000001011011000001;
        10'd483: Q <= 24'b011011000001011011000001;
        10'd484: Q <= 24'b011011000001011011000001;
        10'd485: Q <= 24'b011011000001011011000001;
        10'd486: Q <= 24'b011011000001011011000001;
        10'd487: Q <= 24'b011011000001011011000001;
        10'd488: Q <= 24'b011011000001011011000001;
        10'd489: Q <= 24'b011011000001011011000001;
        10'd490: Q <= 24'b011011000001011011000001;
        10'd491: Q <= 24'b011011000001011011000001;
        10'd492: Q <= 24'b011011000001011011000001;
        10'd493: Q <= 24'b011011000001011011000001;
        10'd494: Q <= 24'b011011000001011011000001;
        10'd495: Q <= 24'b011011000001011011000001;
        10'd496: Q <= 24'b011011000001011011000001;
        10'd497: Q <= 24'b011011000001011011000001;
        10'd498: Q <= 24'b011011000001011011000001;
        10'd499: Q <= 24'b011011000001011011000001;
        10'd500: Q <= 24'b011011000001011011000001;
        10'd501: Q <= 24'b011011000001011011000001;
        10'd502: Q <= 24'b011011000001011011000001;
        10'd503: Q <= 24'b011011000001011011000001;
        10'd504: Q <= 24'b011011000001011011000001;
        10'd505: Q <= 24'b011011000001011011000001;
        10'd506: Q <= 24'b011011000001011011000001;
        10'd507: Q <= 24'b011011000001011011000001;
        10'd508: Q <= 24'b011011000001011011000001;
        10'd509: Q <= 24'b011011000001011011000001;
        10'd510: Q <= 24'b011011000001011011000001;
        10'd511: Q <= 24'b011011000001011011000001;
        10'd512: Q <= 24'b110011011001110011011001;
        10'd513: Q <= 24'b110011011001110011011001;
        10'd514: Q <= 24'b110011011001110011011001;
        10'd515: Q <= 24'b110011011001110011011001;
        10'd516: Q <= 24'b110011011001110011011001;
        10'd517: Q <= 24'b110011011001110011011001;
        10'd518: Q <= 24'b110011011001110011011001;
        10'd519: Q <= 24'b110011011001110011011001;
        10'd520: Q <= 24'b110011011001110011011001;
        10'd521: Q <= 24'b110011011001110011011001;
        10'd522: Q <= 24'b110011011001110011011001;
        10'd523: Q <= 24'b110011011001110011011001;
        10'd524: Q <= 24'b110011011001110011011001;
        10'd525: Q <= 24'b110011011001110011011001;
        10'd526: Q <= 24'b110011011001110011011001;
        10'd527: Q <= 24'b110011011001110011011001;
        10'd528: Q <= 24'b110011011001110011011001;
        10'd529: Q <= 24'b110011011001110011011001;
        10'd530: Q <= 24'b110011011001110011011001;
        10'd531: Q <= 24'b110011011001110011011001;
        10'd532: Q <= 24'b110011011001110011011001;
        10'd533: Q <= 24'b110011011001110011011001;
        10'd534: Q <= 24'b110011011001110011011001;
        10'd535: Q <= 24'b110011011001110011011001;
        10'd536: Q <= 24'b110011011001110011011001;
        10'd537: Q <= 24'b110011011001110011011001;
        10'd538: Q <= 24'b110011011001110011011001;
        10'd539: Q <= 24'b110011011001110011011001;
        10'd540: Q <= 24'b110011011001110011011001;
        10'd541: Q <= 24'b110011011001110011011001;
        10'd542: Q <= 24'b110011011001110011011001;
        10'd543: Q <= 24'b110011011001110011011001;
        10'd544: Q <= 24'b101000010100101000010100;
        10'd545: Q <= 24'b101000010100101000010100;
        10'd546: Q <= 24'b101000010100101000010100;
        10'd547: Q <= 24'b101000010100101000010100;
        10'd548: Q <= 24'b101000010100101000010100;
        10'd549: Q <= 24'b101000010100101000010100;
        10'd550: Q <= 24'b101000010100101000010100;
        10'd551: Q <= 24'b101000010100101000010100;
        10'd552: Q <= 24'b101000010100101000010100;
        10'd553: Q <= 24'b101000010100101000010100;
        10'd554: Q <= 24'b101000010100101000010100;
        10'd555: Q <= 24'b101000010100101000010100;
        10'd556: Q <= 24'b101000010100101000010100;
        10'd557: Q <= 24'b101000010100101000010100;
        10'd558: Q <= 24'b101000010100101000010100;
        10'd559: Q <= 24'b101000010100101000010100;
        10'd560: Q <= 24'b101000010100101000010100;
        10'd561: Q <= 24'b101000010100101000010100;
        10'd562: Q <= 24'b101000010100101000010100;
        10'd563: Q <= 24'b101000010100101000010100;
        10'd564: Q <= 24'b101000010100101000010100;
        10'd565: Q <= 24'b101000010100101000010100;
        10'd566: Q <= 24'b101000010100101000010100;
        10'd567: Q <= 24'b101000010100101000010100;
        10'd568: Q <= 24'b101000010100101000010100;
        10'd569: Q <= 24'b101000010100101000010100;
        10'd570: Q <= 24'b101000010100101000010100;
        10'd571: Q <= 24'b101000010100101000010100;
        10'd572: Q <= 24'b101000010100101000010100;
        10'd573: Q <= 24'b101000010100101000010100;
        10'd574: Q <= 24'b101000010100101000010100;
        10'd575: Q <= 24'b101000010100101000010100;
        10'd576: Q <= 24'b001101010000001101010000;
        10'd577: Q <= 24'b001101010000001101010000;
        10'd578: Q <= 24'b001101010000001101010000;
        10'd579: Q <= 24'b001101010000001101010000;
        10'd580: Q <= 24'b001101010000001101010000;
        10'd581: Q <= 24'b001101010000001101010000;
        10'd582: Q <= 24'b001101010000001101010000;
        10'd583: Q <= 24'b001101010000001101010000;
        10'd584: Q <= 24'b001101010000001101010000;
        10'd585: Q <= 24'b001101010000001101010000;
        10'd586: Q <= 24'b001101010000001101010000;
        10'd587: Q <= 24'b001101010000001101010000;
        10'd588: Q <= 24'b001101010000001101010000;
        10'd589: Q <= 24'b001101010000001101010000;
        10'd590: Q <= 24'b001101010000001101010000;
        10'd591: Q <= 24'b001101010000001101010000;
        10'd592: Q <= 24'b011101101001011101101001;
        10'd593: Q <= 24'b011101101001011101101001;
        10'd594: Q <= 24'b011101101001011101101001;
        10'd595: Q <= 24'b011101101001011101101001;
        10'd596: Q <= 24'b011101101001011101101001;
        10'd597: Q <= 24'b011101101001011101101001;
        10'd598: Q <= 24'b011101101001011101101001;
        10'd599: Q <= 24'b011101101001011101101001;
        10'd600: Q <= 24'b011101101001011101101001;
        10'd601: Q <= 24'b011101101001011101101001;
        10'd602: Q <= 24'b011101101001011101101001;
        10'd603: Q <= 24'b011101101001011101101001;
        10'd604: Q <= 24'b011101101001011101101001;
        10'd605: Q <= 24'b011101101001011101101001;
        10'd606: Q <= 24'b011101101001011101101001;
        10'd607: Q <= 24'b011101101001011101101001;
        10'd608: Q <= 24'b001001110110001001110110;
        10'd609: Q <= 24'b001001110110001001110110;
        10'd610: Q <= 24'b001001110110001001110110;
        10'd611: Q <= 24'b001001110110001001110110;
        10'd612: Q <= 24'b001001110110001001110110;
        10'd613: Q <= 24'b001001110110001001110110;
        10'd614: Q <= 24'b001001110110001001110110;
        10'd615: Q <= 24'b001001110110001001110110;
        10'd616: Q <= 24'b001001110110001001110110;
        10'd617: Q <= 24'b001001110110001001110110;
        10'd618: Q <= 24'b001001110110001001110110;
        10'd619: Q <= 24'b001001110110001001110110;
        10'd620: Q <= 24'b001001110110001001110110;
        10'd621: Q <= 24'b001001110110001001110110;
        10'd622: Q <= 24'b001001110110001001110110;
        10'd623: Q <= 24'b001001110110001001110110;
        10'd624: Q <= 24'b101001010010101001010010;
        10'd625: Q <= 24'b101001010010101001010010;
        10'd626: Q <= 24'b101001010010101001010010;
        10'd627: Q <= 24'b101001010010101001010010;
        10'd628: Q <= 24'b101001010010101001010010;
        10'd629: Q <= 24'b101001010010101001010010;
        10'd630: Q <= 24'b101001010010101001010010;
        10'd631: Q <= 24'b101001010010101001010010;
        10'd632: Q <= 24'b101001010010101001010010;
        10'd633: Q <= 24'b101001010010101001010010;
        10'd634: Q <= 24'b101001010010101001010010;
        10'd635: Q <= 24'b101001010010101001010010;
        10'd636: Q <= 24'b101001010010101001010010;
        10'd637: Q <= 24'b101001010010101001010010;
        10'd638: Q <= 24'b101001010010101001010010;
        10'd639: Q <= 24'b101001010010101001010010;
        10'd640: Q <= 24'b011011010010011011010010;
        10'd641: Q <= 24'b011011010010011011010010;
        10'd642: Q <= 24'b011011010010011011010010;
        10'd643: Q <= 24'b011011010010011011010010;
        10'd644: Q <= 24'b011011010010011011010010;
        10'd645: Q <= 24'b011011010010011011010010;
        10'd646: Q <= 24'b011011010010011011010010;
        10'd647: Q <= 24'b011011010010011011010010;
        10'd648: Q <= 24'b001000111001001000111001;
        10'd649: Q <= 24'b001000111001001000111001;
        10'd650: Q <= 24'b001000111001001000111001;
        10'd651: Q <= 24'b001000111001001000111001;
        10'd652: Q <= 24'b001000111001001000111001;
        10'd653: Q <= 24'b001000111001001000111001;
        10'd654: Q <= 24'b001000111001001000111001;
        10'd655: Q <= 24'b001000111001001000111001;
        10'd656: Q <= 24'b110010111100110010111100;
        10'd657: Q <= 24'b110010111100110010111100;
        10'd658: Q <= 24'b110010111100110010111100;
        10'd659: Q <= 24'b110010111100110010111100;
        10'd660: Q <= 24'b110010111100110010111100;
        10'd661: Q <= 24'b110010111100110010111100;
        10'd662: Q <= 24'b110010111100110010111100;
        10'd663: Q <= 24'b110010111100110010111100;
        10'd664: Q <= 24'b101011100010101011100010;
        10'd665: Q <= 24'b101011100010101011100010;
        10'd666: Q <= 24'b101011100010101011100010;
        10'd667: Q <= 24'b101011100010101011100010;
        10'd668: Q <= 24'b101011100010101011100010;
        10'd669: Q <= 24'b101011100010101011100010;
        10'd670: Q <= 24'b101011100010101011100010;
        10'd671: Q <= 24'b101011100010101011100010;
        10'd672: Q <= 24'b001100011101001100011101;
        10'd673: Q <= 24'b001100011101001100011101;
        10'd674: Q <= 24'b001100011101001100011101;
        10'd675: Q <= 24'b001100011101001100011101;
        10'd676: Q <= 24'b001100011101001100011101;
        10'd677: Q <= 24'b001100011101001100011101;
        10'd678: Q <= 24'b001100011101001100011101;
        10'd679: Q <= 24'b001100011101001100011101;
        10'd680: Q <= 24'b000011000001000011000001;
        10'd681: Q <= 24'b000011000001000011000001;
        10'd682: Q <= 24'b000011000001000011000001;
        10'd683: Q <= 24'b000011000001000011000001;
        10'd684: Q <= 24'b000011000001000011000001;
        10'd685: Q <= 24'b000011000001000011000001;
        10'd686: Q <= 24'b000011000001000011000001;
        10'd687: Q <= 24'b000011000001000011000001;
        10'd688: Q <= 24'b011101111111011101111111;
        10'd689: Q <= 24'b011101111111011101111111;
        10'd690: Q <= 24'b011101111111011101111111;
        10'd691: Q <= 24'b011101111111011101111111;
        10'd692: Q <= 24'b011101111111011101111111;
        10'd693: Q <= 24'b011101111111011101111111;
        10'd694: Q <= 24'b011101111111011101111111;
        10'd695: Q <= 24'b011101111111011101111111;
        10'd696: Q <= 24'b010000100110010000100110;
        10'd697: Q <= 24'b010000100110010000100110;
        10'd698: Q <= 24'b010000100110010000100110;
        10'd699: Q <= 24'b010000100110010000100110;
        10'd700: Q <= 24'b010000100110010000100110;
        10'd701: Q <= 24'b010000100110010000100110;
        10'd702: Q <= 24'b010000100110010000100110;
        10'd703: Q <= 24'b010000100110010000100110;
        10'd704: Q <= 24'b001100110101001100110101;
        10'd705: Q <= 24'b001100110101001100110101;
        10'd706: Q <= 24'b001100110101001100110101;
        10'd707: Q <= 24'b001100110101001100110101;
        10'd708: Q <= 24'b011110110110011110110110;
        10'd709: Q <= 24'b011110110110011110110110;
        10'd710: Q <= 24'b011110110110011110110110;
        10'd711: Q <= 24'b011110110110011110110110;
        10'd712: Q <= 24'b101100111111101100111111;
        10'd713: Q <= 24'b101100111111101100111111;
        10'd714: Q <= 24'b101100111111101100111111;
        10'd715: Q <= 24'b101100111111101100111111;
        10'd716: Q <= 24'b100101011001100101011001;
        10'd717: Q <= 24'b100101011001100101011001;
        10'd718: Q <= 24'b100101011001100101011001;
        10'd719: Q <= 24'b100101011001100101011001;
        10'd720: Q <= 24'b101101000010101101000010;
        10'd721: Q <= 24'b101101000010101101000010;
        10'd722: Q <= 24'b101101000010101101000010;
        10'd723: Q <= 24'b101101000010101101000010;
        10'd724: Q <= 24'b001000010111001000010111;
        10'd725: Q <= 24'b001000010111001000010111;
        10'd726: Q <= 24'b001000010111001000010111;
        10'd727: Q <= 24'b001000010111001000010111;
        10'd728: Q <= 24'b100000101110100000101110;
        10'd729: Q <= 24'b100000101110100000101110;
        10'd730: Q <= 24'b100000101110100000101110;
        10'd731: Q <= 24'b100000101110100000101110;
        10'd732: Q <= 24'b010110010010010110010010;
        10'd733: Q <= 24'b010110010010010110010010;
        10'd734: Q <= 24'b010110010010010110010010;
        10'd735: Q <= 24'b010110010010010110010010;
        10'd736: Q <= 24'b010100110101010100110101;
        10'd737: Q <= 24'b010100110101010100110101;
        10'd738: Q <= 24'b010100110101010100110101;
        10'd739: Q <= 24'b010100110101010100110101;
        10'd740: Q <= 24'b100011000000100011000000;
        10'd741: Q <= 24'b100011000000100011000000;
        10'd742: Q <= 24'b100011000000100011000000;
        10'd743: Q <= 24'b100011000000100011000000;
        10'd744: Q <= 24'b000000111000000000111000;
        10'd745: Q <= 24'b000000111000000000111000;
        10'd746: Q <= 24'b000000111000000000111000;
        10'd747: Q <= 24'b000000111000000000111000;
        10'd748: Q <= 24'b101111100110101111100110;
        10'd749: Q <= 24'b101111100110101111100110;
        10'd750: Q <= 24'b101111100110101111100110;
        10'd751: Q <= 24'b101111100110101111100110;
        10'd752: Q <= 24'b010111000100010111000100;
        10'd753: Q <= 24'b010111000100010111000100;
        10'd754: Q <= 24'b010111000100010111000100;
        10'd755: Q <= 24'b010111000100010111000100;
        10'd756: Q <= 24'b010100111011010100111011;
        10'd757: Q <= 24'b010100111011010100111011;
        10'd758: Q <= 24'b010100111011010100111011;
        10'd759: Q <= 24'b010100111011010100111011;
        10'd760: Q <= 24'b100110001111100110001111;
        10'd761: Q <= 24'b100110001111100110001111;
        10'd762: Q <= 24'b100110001111100110001111;
        10'd763: Q <= 24'b100110001111100110001111;
        10'd764: Q <= 24'b000100101000000100101000;
        10'd765: Q <= 24'b000100101000000100101000;
        10'd766: Q <= 24'b000100101000000100101000;
        10'd767: Q <= 24'b000100101000000100101000;
        10'd768: Q <= 24'b001110001110001110001110;
        10'd769: Q <= 24'b001110001110001110001110;
        10'd770: Q <= 24'b010011001011010011001011;
        10'd771: Q <= 24'b010011001011010011001011;
        10'd772: Q <= 24'b110000100110110000100110;
        10'd773: Q <= 24'b110000100110110000100110;
        10'd774: Q <= 24'b100110101010100110101010;
        10'd775: Q <= 24'b100110101010100110101010;
        10'd776: Q <= 24'b001010001000001010001000;
        10'd777: Q <= 24'b001010001000001010001000;
        10'd778: Q <= 24'b010111001001010111001001;
        10'd779: Q <= 24'b010111001001010111001001;
        10'd780: Q <= 24'b101000111001101000111001;
        10'd781: Q <= 24'b101000111001101000111001;
        10'd782: Q <= 24'b101001010111101001010111;
        10'd783: Q <= 24'b101001010111101001010111;
        10'd784: Q <= 24'b100101100010100101100010;
        10'd785: Q <= 24'b100101100010100101100010;
        10'd786: Q <= 24'b010111111110010111111110;
        10'd787: Q <= 24'b010111111110010111111110;
        10'd788: Q <= 24'b101100110100101100110100;
        10'd789: Q <= 24'b101100110100101100110100;
        10'd790: Q <= 24'b010110011110010110011110;
        10'd791: Q <= 24'b010110011110010110011110;
        10'd792: Q <= 24'b000111000100000111000100;
        10'd793: Q <= 24'b000111000100000111000100;
        10'd794: Q <= 24'b001100100111001100100111;
        10'd795: Q <= 24'b001100100111001100100111;
        10'd796: Q <= 24'b010110011011010110011011;
        10'd797: Q <= 24'b010110011011010110011011;
        10'd798: Q <= 24'b100100001111100100001111;
        10'd799: Q <= 24'b100100001111100100001111;
        10'd800: Q <= 24'b011101111011011101111011;
        10'd801: Q <= 24'b011101111011011101111011;
        10'd802: Q <= 24'b010100101000010100101000;
        10'd803: Q <= 24'b010100101000010100101000;
        10'd804: Q <= 24'b000000100001000000100001;
        10'd805: Q <= 24'b000000100001000000100001;
        10'd806: Q <= 24'b101100110001101100110001;
        10'd807: Q <= 24'b101100110001101100110001;
        10'd808: Q <= 24'b001001111000001001111000;
        10'd809: Q <= 24'b001001111000001001111000;
        10'd810: Q <= 24'b100111010001100111010001;
        10'd811: Q <= 24'b100111010001100111010001;
        10'd812: Q <= 24'b011110111001011110111001;
        10'd813: Q <= 24'b011110111001011110111001;
        10'd814: Q <= 24'b001010001010001010001010;
        10'd815: Q <= 24'b001010001010001010001010;
        10'd816: Q <= 24'b100000000111100000000111;
        10'd817: Q <= 24'b100000000111100000000111;
        10'd818: Q <= 24'b100011100101100011100101;
        10'd819: Q <= 24'b100011100101100011100101;
        10'd820: Q <= 24'b100100000000100100000000;
        10'd821: Q <= 24'b100100000000100100000000;
        10'd822: Q <= 24'b010010101101010010101101;
        10'd823: Q <= 24'b010010101101010010101101;
        10'd824: Q <= 24'b011011011100011011011100;
        10'd825: Q <= 24'b011011011100011011011100;
        10'd826: Q <= 24'b110010110101110010110101;
        10'd827: Q <= 24'b110010110101110010110101;
        10'd828: Q <= 24'b000101001011000101001011;
        10'd829: Q <= 24'b000101001011000101001011;
        10'd830: Q <= 24'b000100100001000100100001;
        10'd831: Q <= 24'b000100100001000100100001;
        10'd832: Q <= 24'b100001101010100001101010;
        10'd833: Q <= 24'b001101110101001101110101;
        10'd834: Q <= 24'b101101110111101101110111;
        10'd835: Q <= 24'b100000111110100000111110;
        10'd836: Q <= 24'b010000000101010000000101;
        10'd837: Q <= 24'b011101010010011101010010;
        10'd838: Q <= 24'b010010111100010010111100;
        10'd839: Q <= 24'b011010111010011010111010;
        10'd840: Q <= 24'b001101110110001101110110;
        10'd841: Q <= 24'b101011010111101011010111;
        10'd842: Q <= 24'b100001100110100001100110;
        10'd843: Q <= 24'b010001110111010001110111;
        10'd844: Q <= 24'b010000000010010000000010;
        10'd845: Q <= 24'b000110010011000110010011;
        10'd846: Q <= 24'b010001000100010001000100;
        10'd847: Q <= 24'b101011110100101011110100;
        10'd848: Q <= 24'b101000100010101000100010;
        10'd849: Q <= 24'b100110100010100110100010;
        10'd850: Q <= 24'b001000110001001000110001;
        10'd851: Q <= 24'b100000110011100000110011;
        10'd852: Q <= 24'b001011110101001011110101;
        10'd853: Q <= 24'b101011010101101011010101;
        10'd854: Q <= 24'b000100111111000100111111;
        10'd855: Q <= 24'b010000100111010000100111;
        10'd856: Q <= 24'b011001101101011001101101;
        10'd857: Q <= 24'b100000101010100000101010;
        10'd858: Q <= 24'b100111110101100111110101;
        10'd859: Q <= 24'b000101110111000101110111;
        10'd860: Q <= 24'b110010010100110010010100;
        10'd861: Q <= 24'b011111110101011111110101;
        10'd862: Q <= 24'b100011111010100011111010;
        10'd863: Q <= 24'b011000110000011000110000;
        10'd864: Q <= 24'b001010000001001010000001;
        10'd865: Q <= 24'b000100001100000100001100;
        10'd866: Q <= 24'b100100100001100100100001;
        10'd867: Q <= 24'b001011011101001011011101;
        10'd868: Q <= 24'b100101010100100101010100;
        10'd869: Q <= 24'b100110000101100110000101;
        10'd870: Q <= 24'b100100000100100100000100;
        10'd871: Q <= 24'b001110101011001110101011;
        10'd872: Q <= 24'b101001111111101001111111;
        10'd873: Q <= 24'b010110110101010110110101;
        10'd874: Q <= 24'b001110111000001110111000;
        10'd875: Q <= 24'b011100110111011100110111;
        10'd876: Q <= 24'b011011111101011011111101;
        10'd877: Q <= 24'b101011100101101011100101;
        10'd878: Q <= 24'b011001110011011001110011;
        10'd879: Q <= 24'b011010100111011010100111;
        10'd880: Q <= 24'b101111101010101111101010;
        10'd881: Q <= 24'b101111000111101111000111;
        10'd882: Q <= 24'b100001101100100001101100;
        10'd883: Q <= 24'b001011110100001011110100;
        10'd884: Q <= 24'b000011101001000011101001;
        10'd885: Q <= 24'b110011010001110011010001;
        10'd886: Q <= 24'b101001100110101001100110;
        10'd887: Q <= 24'b010110000001010110000001;
        10'd888: Q <= 24'b010001001100010001001100;
        10'd889: Q <= 24'b100011110000100011110000;
        10'd890: Q <= 24'b001011010011001011010011;
        10'd891: Q <= 24'b011001100101011001100101;
        10'd892: Q <= 24'b101001011001101001011001;
        10'd893: Q <= 24'b001001000111001001000111;
        10'd894: Q <= 24'b101011001001101011001001;
        10'd895: Q <= 24'b000000010001000000010001;
        10'd896: Q <= 24'b000000000000000000010001;
        10'd897: Q <= 24'b000000000000110011110000;
        10'd898: Q <= 24'b000000000000101011001001;
        10'd899: Q <= 24'b000000000000001000111000;
        10'd900: Q <= 24'b000000000000001001000111;
        10'd901: Q <= 24'b000000000000101010111010;
        10'd902: Q <= 24'b000000000000101001011001;
        10'd903: Q <= 24'b000000000000001010101000;
        10'd904: Q <= 24'b000000000000011001100101;
        10'd905: Q <= 24'b000000000000011010011100;
        10'd906: Q <= 24'b000000000000001011010011;
        10'd907: Q <= 24'b000000000000101000101110;
        10'd908: Q <= 24'b000000000000100011110000;
        10'd909: Q <= 24'b000000000000010000010001;
        10'd910: Q <= 24'b000000000000010001001100;
        10'd911: Q <= 24'b000000000000100010110101;
        10'd912: Q <= 24'b000000000000010110000001;
        10'd913: Q <= 24'b000000000000011110000000;
        10'd914: Q <= 24'b000000000000101001100110;
        10'd915: Q <= 24'b000000000000001010011011;
        10'd916: Q <= 24'b000000000000110011010001;
        10'd917: Q <= 24'b000000000000000000110000;
        10'd918: Q <= 24'b000000000000000011101001;
        10'd919: Q <= 24'b000000000000110000011000;
        10'd920: Q <= 24'b000000000000001011110100;
        10'd921: Q <= 24'b000000000000101000001101;
        10'd922: Q <= 24'b000000000000100001101100;
        10'd923: Q <= 24'b000000000000010010010101;
        10'd924: Q <= 24'b000000000000101111000111;
        10'd925: Q <= 24'b000000000000000100111010;
        10'd926: Q <= 24'b000000000000101111101010;
        10'd927: Q <= 24'b000000000000000100010111;
        10'd928: Q <= 24'b000000000000011010100111;
        10'd929: Q <= 24'b000000000000011001011010;
        10'd930: Q <= 24'b000000000000011001110011;
        10'd931: Q <= 24'b000000000000011010001110;
        10'd932: Q <= 24'b000000000000101011100101;
        10'd933: Q <= 24'b000000000000001000011100;
        10'd934: Q <= 24'b000000000000011011111101;
        10'd935: Q <= 24'b000000000000011000000100;
        10'd936: Q <= 24'b000000000000011100110111;
        10'd937: Q <= 24'b000000000000010111001010;
        10'd938: Q <= 24'b000000000000001110111000;
        10'd939: Q <= 24'b000000000000100101001001;
        10'd940: Q <= 24'b000000000000010110110101;
        10'd941: Q <= 24'b000000000000011101001100;
        10'd942: Q <= 24'b000000000000101001111111;
        10'd943: Q <= 24'b000000000000001010000010;
        10'd944: Q <= 24'b000000000000001110101011;
        10'd945: Q <= 24'b000000000000100101010110;
        10'd946: Q <= 24'b000000000000100100000100;
        10'd947: Q <= 24'b000000000000001111111101;
        10'd948: Q <= 24'b000000000000100110000101;
        10'd949: Q <= 24'b000000000000001101111100;
        10'd950: Q <= 24'b000000000000100101010100;
        10'd951: Q <= 24'b000000000000001110101101;
        10'd952: Q <= 24'b000000000000001011011101;
        10'd953: Q <= 24'b000000000000101000100100;
        10'd954: Q <= 24'b000000000000100100100001;
        10'd955: Q <= 24'b000000000000001111100000;
        10'd956: Q <= 24'b000000000000000100001100;
        10'd957: Q <= 24'b000000000000101111110101;
        10'd958: Q <= 24'b000000000000001010000001;
        10'd959: Q <= 24'b000000000000101010000000;
        10'd960: Q <= 24'b000000000000011000110000;
        10'd961: Q <= 24'b000000000000011011010001;
        10'd962: Q <= 24'b000000000000100011111010;
        10'd963: Q <= 24'b000000000000010000000111;
        10'd964: Q <= 24'b000000000000011111110101;
        10'd965: Q <= 24'b000000000000010100001100;
        10'd966: Q <= 24'b000000000000110010010100;
        10'd967: Q <= 24'b000000000000000001101101;
        10'd968: Q <= 24'b000000000000000101110111;
        10'd969: Q <= 24'b000000000000101110001010;
        10'd970: Q <= 24'b000000000000100111110101;
        10'd971: Q <= 24'b000000000000001100001100;
        10'd972: Q <= 24'b000000000000100000101010;
        10'd973: Q <= 24'b000000000000010011010111;
        10'd974: Q <= 24'b000000000000011001101101;
        10'd975: Q <= 24'b000000000000011010010100;
        10'd976: Q <= 24'b000000000000010000100111;
        10'd977: Q <= 24'b000000000000100011011010;
        10'd978: Q <= 24'b000000000000000100111111;
        10'd979: Q <= 24'b000000000000101111000010;
        10'd980: Q <= 24'b000000000000101011010101;
        10'd981: Q <= 24'b000000000000001000101100;
        10'd982: Q <= 24'b000000000000001011110101;
        10'd983: Q <= 24'b000000000000101000001100;
        10'd984: Q <= 24'b000000000000100000110011;
        10'd985: Q <= 24'b000000000000010011001110;
        10'd986: Q <= 24'b000000000000001000110001;
        10'd987: Q <= 24'b000000000000101011010000;
        10'd988: Q <= 24'b000000000000100110100010;
        10'd989: Q <= 24'b000000000000001101011111;
        10'd990: Q <= 24'b000000000000101000100010;
        10'd991: Q <= 24'b000000000000001011011111;
        10'd992: Q <= 24'b000000000000101011110100;
        10'd993: Q <= 24'b000000000000001000001101;
        10'd994: Q <= 24'b000000000000010001000100;
        10'd995: Q <= 24'b000000000000100010111101;
        10'd996: Q <= 24'b000000000000000110010011;
        10'd997: Q <= 24'b000000000000101101101110;
        10'd998: Q <= 24'b000000000000010000000010;
        10'd999: Q <= 24'b000000000000100011111111;
        10'd1000: Q <=24'b000000000000010001110111;
        10'd1001: Q <=24'b000000000000100010001010;
        10'd1002: Q <=24'b000000000000100001100110;
        10'd1003: Q <=24'b000000000000010010011011;
        10'd1004: Q <=24'b000000000000101011010111;
        10'd1005: Q <=24'b000000000000001000101010;
        10'd1006: Q <=24'b000000000000001101110110;
        10'd1007: Q <=24'b000000000000100110001011;
        10'd1008: Q <=24'b000000000000011010111010;
        10'd1009: Q <=24'b000000000000011001000111;
        10'd1010: Q <=24'b000000000000010010111100;
        10'd1011: Q <=24'b000000000000100001000101;
        10'd1012: Q <=24'b000000000000011101010010;
        10'd1013: Q <=24'b000000000000010110101111;
        10'd1014: Q <=24'b000000000000010000000101;
        10'd1015: Q <=24'b000000000000100011111100;
        10'd1016: Q <=24'b000000000000100000111110;
        10'd1017: Q <=24'b000000000000010011000011;
        10'd1018: Q <=24'b000000000000101101110111;
        10'd1019: Q <=24'b000000000000000110001010;
        10'd1020: Q <=24'b000000000000001101110101;
        10'd1021: Q <=24'b000000000000100110001100;
        10'd1022: Q <=24'b000000000000100001101010;
        10'd1023: Q <=24'b000000000000010010010111;
        endcase end         
        end
`elsif OP1
    always@(posedge clk)
        begin
        if(REN == 1'b1) begin
        case(A)
        9'd0:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd1:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd2:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd3:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd4:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd5:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd6:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd7:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd8:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd9:   Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd10:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd11:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd12:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd13:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd14:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd15:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd16:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd17:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd18:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd19:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd20:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd21:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd22:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd23:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd24:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd25:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd26:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd27:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd28:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd29:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd30:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd31:  Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd32:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd33:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd34:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd35:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd36:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd37:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd38:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd39:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd40:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd41:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd42:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd43:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd44:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd45:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd46:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd47:  Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd48:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd49:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd50:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd51:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd52:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd53:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd54:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd55:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd56:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd57:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd58:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd59:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd60:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd61:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd62:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd63:  Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd64:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd65:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd66:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd67:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd68:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd69:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd70:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd71:  Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd72:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd73:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd74:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd75:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd76:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd77:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd78:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd79:  Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd80:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd81:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd82:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd83:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd84:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd85:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd86:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd87:  Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd88:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd89:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd90:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd91:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd92:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd93:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd94:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd95:  Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd96:  Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd97:  Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd98:  Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd99:  Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd100: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd101: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd102: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd103: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd104: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd105: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd106: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd107: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd108: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd109: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd110: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd111: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd112: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd113: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd114: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd115: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd116: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd117: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd118: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd119: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd120: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd121: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd122: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd123: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd124: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd125: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd126: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd127: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd128: Q <= 48'b000100101000000100101000000100101000000100101000;
        9'd129: Q <= 48'b000100101000000100101000000100101000000100101000;
        9'd130: Q <= 48'b100110001111100110001111100110001111100110001111;
        9'd131: Q <= 48'b100110001111100110001111100110001111100110001111;
        9'd132: Q <= 48'b010100111011010100111011010100111011010100111011;
        9'd133: Q <= 48'b010100111011010100111011010100111011010100111011;
        9'd134: Q <= 48'b010111000100010111000100010111000100010111000100;
        9'd135: Q <= 48'b010111000100010111000100010111000100010111000100;
        9'd136: Q <= 48'b101111100110101111100110101111100110101111100110;
        9'd137: Q <= 48'b101111100110101111100110101111100110101111100110;
        9'd138: Q <= 48'b000000111000000000111000000000111000000000111000;
        9'd139: Q <= 48'b000000111000000000111000000000111000000000111000;
        9'd140: Q <= 48'b100011000000100011000000100011000000100011000000;
        9'd141: Q <= 48'b100011000000100011000000100011000000100011000000;
        9'd142: Q <= 48'b010100110101010100110101010100110101010100110101;
        9'd143: Q <= 48'b010100110101010100110101010100110101010100110101;
        9'd144: Q <= 48'b010110010010010110010010010110010010010110010010;
        9'd145: Q <= 48'b010110010010010110010010010110010010010110010010;
        9'd146: Q <= 48'b100000101110100000101110100000101110100000101110;
        9'd147: Q <= 48'b100000101110100000101110100000101110100000101110;
        9'd148: Q <= 48'b001000010111001000010111001000010111001000010111;
        9'd149: Q <= 48'b001000010111001000010111001000010111001000010111;
        9'd150: Q <= 48'b101101000010101101000010101101000010101101000010;
        9'd151: Q <= 48'b101101000010101101000010101101000010101101000010;
        9'd152: Q <= 48'b100101011001100101011001100101011001100101011001;
        9'd153: Q <= 48'b100101011001100101011001100101011001100101011001;
        9'd154: Q <= 48'b101100111111101100111111101100111111101100111111;
        9'd155: Q <= 48'b101100111111101100111111101100111111101100111111;
        9'd156: Q <= 48'b011110110110011110110110011110110110011110110110;
        9'd157: Q <= 48'b011110110110011110110110011110110110011110110110;
        9'd158: Q <= 48'b001100110101001100110101001100110101001100110101;
        9'd159: Q <= 48'b001100110101001100110101001100110101001100110101;
        9'd160: Q <= 48'b000100100001000100100001000100100001000100100001;
        9'd161: Q <= 48'b000101001011000101001011000101001011000101001011;
        9'd162: Q <= 48'b110010110101110010110101110010110101110010110101;
        9'd163: Q <= 48'b011011011100011011011100011011011100011011011100;
        9'd164: Q <= 48'b010010101101010010101101010010101101010010101101;
        9'd165: Q <= 48'b100100000000100100000000100100000000100100000000;
        9'd166: Q <= 48'b100011100101100011100101100011100101100011100101;
        9'd167: Q <= 48'b100000000111100000000111100000000111100000000111;
        9'd168: Q <= 48'b001010001010001010001010001010001010001010001010;
        9'd169: Q <= 48'b011110111001011110111001011110111001011110111001;
        9'd170: Q <= 48'b100111010001100111010001100111010001100111010001;
        9'd171: Q <= 48'b001001111000001001111000001001111000001001111000;
        9'd172: Q <= 48'b101100110001101100110001101100110001101100110001;
        9'd173: Q <= 48'b000000100001000000100001000000100001000000100001;
        9'd174: Q <= 48'b010100101000010100101000010100101000010100101000;
        9'd175: Q <= 48'b011101111011011101111011011101111011011101111011;
        9'd176: Q <= 48'b100100001111100100001111100100001111100100001111;
        9'd177: Q <= 48'b010110011011010110011011010110011011010110011011;
        9'd178: Q <= 48'b001100100111001100100111001100100111001100100111;
        9'd179: Q <= 48'b000111000100000111000100000111000100000111000100;
        9'd180: Q <= 48'b010110011110010110011110010110011110010110011110;
        9'd181: Q <= 48'b101100110100101100110100101100110100101100110100;
        9'd182: Q <= 48'b010111111110010111111110010111111110010111111110;
        9'd183: Q <= 48'b100101100010100101100010100101100010100101100010;
        9'd184: Q <= 48'b101001010111101001010111101001010111101001010111;
        9'd185: Q <= 48'b101000111001101000111001101000111001101000111001;
        9'd186: Q <= 48'b010111001001010111001001010111001001010111001001;
        9'd187: Q <= 48'b001010001000001010001000001010001000001010001000;
        9'd188: Q <= 48'b100110101010100110101010100110101010100110101010;
        9'd189: Q <= 48'b110000100110110000100110110000100110110000100110;
        9'd190: Q <= 48'b010011001011010011001011010011001011010011001011;
        9'd191: Q <= 48'b001110001110001110001110001110001110001110001110;
        9'd192: Q <= 48'b000000010001000000010001101011001001101011001001;
        9'd193: Q <= 48'b001001000111001001000111101001011001101001011001;
        9'd194: Q <= 48'b011001100101011001100101001011010011001011010011;
        9'd195: Q <= 48'b100011110000100011110000010001001100010001001100;
        9'd196: Q <= 48'b010110000001010110000001101001100110101001100110;
        9'd197: Q <= 48'b110011010001110011010001000011101001000011101001;
        9'd198: Q <= 48'b001011110100001011110100100001101100100001101100;
        9'd199: Q <= 48'b101111000111101111000111101111101010101111101010;
        9'd200: Q <= 48'b011010100111011010100111011001110011011001110011;
        9'd201: Q <= 48'b101011100101101011100101011011111101011011111101;
        9'd202: Q <= 48'b011100110111011100110111001110111000001110111000;
        9'd203: Q <= 48'b010110110101010110110101101001111111101001111111;
        9'd204: Q <= 48'b001110101011001110101011100100000100100100000100;
        9'd205: Q <= 48'b100110000101100110000101100101010100100101010100;
        9'd206: Q <= 48'b001011011101001011011101100100100001100100100001;
        9'd207: Q <= 48'b000100001100000100001100001010000001001010000001;
        9'd208: Q <= 48'b011000110000011000110000100011111010100011111010;
        9'd209: Q <= 48'b011111110101011111110101110010010100110010010100;
        9'd210: Q <= 48'b000101110111000101110111100111110101100111110101;
        9'd211: Q <= 48'b100000101010100000101010011001101101011001101101;
        9'd212: Q <= 48'b010000100111010000100111000100111111000100111111;
        9'd213: Q <= 48'b101011010101101011010101001011110101001011110101;
        9'd214: Q <= 48'b100000110011100000110011001000110001001000110001;
        9'd215: Q <= 48'b100110100010100110100010101000100010101000100010;
        9'd216: Q <= 48'b101011110100101011110100010001000100010001000100;
        9'd217: Q <= 48'b000110010011000110010011010000000010010000000010;
        9'd218: Q <= 48'b010001110111010001110111100001100110100001100110;
        9'd219: Q <= 48'b101011010111101011010111001101110110001101110110;
        9'd220: Q <= 48'b011010111010011010111010010010111100010010111100;
        9'd221: Q <= 48'b011101010010011101010010010000000101010000000101;
        9'd222: Q <= 48'b100000111110100000111110101101110111101101110111;
        9'd223: Q <= 48'b001101110101001101110101100001101010100001101010;
        9'd224: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd225: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd226: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd227: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd228: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd229: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd230: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd231: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd232: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd233: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd234: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd235: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd236: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd237: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd238: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd239: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd240: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd241: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd242: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd243: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd244: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd245: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd246: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd247: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd248: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd249: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd250: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd251: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd252: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd253: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd254: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd255: Q <= 48'b011011000001011011000001011011000001011011000001;
        9'd256: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd257: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd258: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd259: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd260: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd261: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd262: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd263: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd264: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd265: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd266: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd267: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd268: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd269: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd270: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd271: Q <= 48'b110011011001110011011001110011011001110011011001;
        9'd272: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd273: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd274: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd275: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd276: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd277: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd278: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd279: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd280: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd281: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd282: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd283: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd284: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd285: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd286: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd287: Q <= 48'b101000010100101000010100101000010100101000010100;
        9'd288: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd289: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd290: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd291: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd292: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd293: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd294: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd295: Q <= 48'b001101010000001101010000001101010000001101010000;
        9'd296: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd297: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd298: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd299: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd300: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd301: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd302: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd303: Q <= 48'b011101101001011101101001011101101001011101101001;
        9'd304: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd305: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd306: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd307: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd308: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd309: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd310: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd311: Q <= 48'b001001110110001001110110001001110110001001110110;
        9'd312: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd313: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd314: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd315: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd316: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd317: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd318: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd319: Q <= 48'b101001010010101001010010101001010010101001010010;
        9'd320: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd321: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd322: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd323: Q <= 48'b011011010010011011010010011011010010011011010010;
        9'd324: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd325: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd326: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd327: Q <= 48'b001000111001001000111001001000111001001000111001;
        9'd328: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd329: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd330: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd331: Q <= 48'b110010111100110010111100110010111100110010111100;
        9'd332: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd333: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd334: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd335: Q <= 48'b101011100010101011100010101011100010101011100010;
        9'd336: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd337: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd338: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd339: Q <= 48'b001100011101001100011101001100011101001100011101;
        9'd340: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd341: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd342: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd343: Q <= 48'b000011000001000011000001000011000001000011000001;
        9'd344: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd345: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd346: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd347: Q <= 48'b011101111111011101111111011101111111011101111111;
        9'd348: Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd349: Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd350: Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd351: Q <= 48'b010000100110010000100110010000100110010000100110;
        9'd352: Q <= 48'b001100110101001100110101001100110101001100110101;
        9'd353: Q <= 48'b001100110101001100110101001100110101001100110101;
        9'd354: Q <= 48'b011110110110011110110110011110110110011110110110;
        9'd355: Q <= 48'b011110110110011110110110011110110110011110110110;
        9'd356: Q <= 48'b101100111111101100111111101100111111101100111111;
        9'd357: Q <= 48'b101100111111101100111111101100111111101100111111;
        9'd358: Q <= 48'b100101011001100101011001100101011001100101011001;
        9'd359: Q <= 48'b100101011001100101011001100101011001100101011001;
        9'd360: Q <= 48'b101101000010101101000010101101000010101101000010;
        9'd361: Q <= 48'b101101000010101101000010101101000010101101000010;
        9'd362: Q <= 48'b001000010111001000010111001000010111001000010111;
        9'd363: Q <= 48'b001000010111001000010111001000010111001000010111;
        9'd364: Q <= 48'b100000101110100000101110100000101110100000101110;
        9'd365: Q <= 48'b100000101110100000101110100000101110100000101110;
        9'd366: Q <= 48'b010110010010010110010010010110010010010110010010;
        9'd367: Q <= 48'b010110010010010110010010010110010010010110010010;
        9'd368: Q <= 48'b010100110101010100110101010100110101010100110101;
        9'd369: Q <= 48'b010100110101010100110101010100110101010100110101;
        9'd370: Q <= 48'b100011000000100011000000100011000000100011000000;
        9'd371: Q <= 48'b100011000000100011000000100011000000100011000000;
        9'd372: Q <= 48'b000000111000000000111000000000111000000000111000;
        9'd373: Q <= 48'b000000111000000000111000000000111000000000111000;
        9'd374: Q <= 48'b101111100110101111100110101111100110101111100110;
        9'd375: Q <= 48'b101111100110101111100110101111100110101111100110;
        9'd376: Q <= 48'b010111000100010111000100010111000100010111000100;
        9'd377: Q <= 48'b010111000100010111000100010111000100010111000100;
        9'd378: Q <= 48'b010100111011010100111011010100111011010100111011;
        9'd379: Q <= 48'b010100111011010100111011010100111011010100111011;
        9'd380: Q <= 48'b100110001111100110001111100110001111100110001111;
        9'd381: Q <= 48'b100110001111100110001111100110001111100110001111;
        9'd382: Q <= 48'b000100101000000100101000000100101000000100101000;
        9'd383: Q <= 48'b000100101000000100101000000100101000000100101000;
        9'd384: Q <= 48'b001110001110001110001110001110001110001110001110;
        9'd385: Q <= 48'b010011001011010011001011010011001011010011001011;
        9'd386: Q <= 48'b110000100110110000100110110000100110110000100110;
        9'd387: Q <= 48'b100110101010100110101010100110101010100110101010;
        9'd388: Q <= 48'b001010001000001010001000001010001000001010001000;
        9'd389: Q <= 48'b010111001001010111001001010111001001010111001001;
        9'd390: Q <= 48'b101000111001101000111001101000111001101000111001;
        9'd391: Q <= 48'b101001010111101001010111101001010111101001010111;
        9'd392: Q <= 48'b100101100010100101100010100101100010100101100010;
        9'd393: Q <= 48'b010111111110010111111110010111111110010111111110;
        9'd394: Q <= 48'b101100110100101100110100101100110100101100110100;
        9'd395: Q <= 48'b010110011110010110011110010110011110010110011110;
        9'd396: Q <= 48'b000111000100000111000100000111000100000111000100;
        9'd397: Q <= 48'b001100100111001100100111001100100111001100100111;
        9'd398: Q <= 48'b010110011011010110011011010110011011010110011011;
        9'd399: Q <= 48'b100100001111100100001111100100001111100100001111;
        9'd400: Q <= 48'b011101111011011101111011011101111011011101111011;
        9'd401: Q <= 48'b010100101000010100101000010100101000010100101000;
        9'd402: Q <= 48'b000000100001000000100001000000100001000000100001;
        9'd403: Q <= 48'b101100110001101100110001101100110001101100110001;
        9'd404: Q <= 48'b001001111000001001111000001001111000001001111000;
        9'd405: Q <= 48'b100111010001100111010001100111010001100111010001;
        9'd406: Q <= 48'b011110111001011110111001011110111001011110111001;
        9'd407: Q <= 48'b001010001010001010001010001010001010001010001010;
        9'd408: Q <= 48'b100000000111100000000111100000000111100000000111;
        9'd409: Q <= 48'b100011100101100011100101100011100101100011100101;
        9'd410: Q <= 48'b100100000000100100000000100100000000100100000000;
        9'd411: Q <= 48'b010010101101010010101101010010101101010010101101;
        9'd412: Q <= 48'b011011011100011011011100011011011100011011011100;
        9'd413: Q <= 48'b110010110101110010110101110010110101110010110101;
        9'd414: Q <= 48'b000101001011000101001011000101001011000101001011;
        9'd415: Q <= 48'b000100100001000100100001000100100001000100100001;
        9'd416: Q <= 48'b100001101010100001101010001101110101001101110101;
        9'd417: Q <= 48'b101101110111101101110111100000111110100000111110;
        9'd418: Q <= 48'b010000000101010000000101011101010010011101010010;
        9'd419: Q <= 48'b010010111100010010111100011010111010011010111010;
        9'd420: Q <= 48'b001101110110001101110110101011010111101011010111;
        9'd421: Q <= 48'b100001100110100001100110010001110111010001110111;
        9'd422: Q <= 48'b010000000010010000000010000110010011000110010011;
        9'd423: Q <= 48'b010001000100010001000100101011110100101011110100;
        9'd424: Q <= 48'b101000100010101000100010100110100010100110100010;
        9'd425: Q <= 48'b001000110001001000110001100000110011100000110011;
        9'd426: Q <= 48'b001011110101001011110101101011010101101011010101;
        9'd427: Q <= 48'b000100111111000100111111010000100111010000100111;
        9'd428: Q <= 48'b011001101101011001101101100000101010100000101010;
        9'd429: Q <= 48'b100111110101100111110101000101110111000101110111;
        9'd430: Q <= 48'b110010010100110010010100011111110101011111110101;
        9'd431: Q <= 48'b100011111010100011111010011000110000011000110000;
        9'd432: Q <= 48'b001010000001001010000001000100001100000100001100;
        9'd433: Q <= 48'b100100100001100100100001001011011101001011011101;
        9'd434: Q <= 48'b100101010100100101010100100110000101100110000101;
        9'd435: Q <= 48'b100100000100100100000100001110101011001110101011;
        9'd436: Q <= 48'b101001111111101001111111010110110101010110110101;
        9'd437: Q <= 48'b001110111000001110111000011100110111011100110111;
        9'd438: Q <= 48'b011011111101011011111101101011100101101011100101;
        9'd439: Q <= 48'b011001110011011001110011011010100111011010100111;
        9'd440: Q <= 48'b101111101010101111101010101111000111101111000111;
        9'd441: Q <= 48'b100001101100100001101100001011110100001011110100;
        9'd442: Q <= 48'b000011101001000011101001110011010001110011010001;
        9'd443: Q <= 48'b101001100110101001100110010110000001010110000001;
        9'd444: Q <= 48'b010001001100010001001100100011110000100011110000;
        9'd445: Q <= 48'b001011010011001011010011011001100101011001100101;
        9'd446: Q <= 48'b101001011001101001011001001001000111001001000111;
        9'd447: Q <= 48'b101011001001101011001001000000010001000000010001;
        9'd448: Q <= 48'b000000000000000000010001000000000000110011110000;
        9'd449: Q <= 48'b000000000000101011001001000000000000001000111000;
        9'd450: Q <= 48'b000000000000001001000111000000000000101010111010;
        9'd451: Q <= 48'b000000000000101001011001000000000000001010101000;
        9'd452: Q <= 48'b000000000000011001100101000000000000011010011100;
        9'd453: Q <= 48'b000000000000001011010011000000000000101000101110;
        9'd454: Q <= 48'b000000000000100011110000000000000000010000010001;
        9'd455: Q <= 48'b000000000000010001001100000000000000100010110101;
        9'd456: Q <= 48'b000000000000010110000001000000000000011110000000;
        9'd457: Q <= 48'b000000000000101001100110000000000000001010011011;
        9'd458: Q <= 48'b000000000000110011010001000000000000000000110000;
        9'd459: Q <= 48'b000000000000000011101001000000000000110000011000;
        9'd460: Q <= 48'b000000000000001011110100000000000000101000001101;
        9'd461: Q <= 48'b000000000000100001101100000000000000010010010101;
        9'd462: Q <= 48'b000000000000101111000111000000000000000100111010;
        9'd463: Q <= 48'b000000000000101111101010000000000000000100010111;
        9'd464: Q <= 48'b000000000000011010100111000000000000011001011010;
        9'd465: Q <= 48'b000000000000011001110011000000000000011010001110;
        9'd466: Q <= 48'b000000000000101011100101000000000000001000011100;
        9'd467: Q <= 48'b000000000000011011111101000000000000011000000100;
        9'd468: Q <= 48'b000000000000011100110111000000000000010111001010;
        9'd469: Q <= 48'b000000000000001110111000000000000000100101001001;
        9'd470: Q <= 48'b000000000000010110110101000000000000011101001100;
        9'd471: Q <= 48'b000000000000101001111111000000000000001010000010;
        9'd472: Q <= 48'b000000000000001110101011000000000000100101010110;
        9'd473: Q <= 48'b000000000000100100000100000000000000001111111101;
        9'd474: Q <= 48'b000000000000100110000101000000000000001101111100;
        9'd475: Q <= 48'b000000000000100101010100000000000000001110101101;
        9'd476: Q <= 48'b000000000000001011011101000000000000101000100100;
        9'd477: Q <= 48'b000000000000100100100001000000000000001111100000;
        9'd478: Q <= 48'b000000000000000100001100000000000000101111110101;
        9'd479: Q <= 48'b000000000000001010000001000000000000101010000000;
        9'd480: Q <= 48'b000000000000011000110000000000000000011011010001;
        9'd481: Q <= 48'b000000000000100011111010000000000000010000000111;
        9'd482: Q <= 48'b000000000000011111110101000000000000010100001100;
        9'd483: Q <= 48'b000000000000110010010100000000000000000001101101;
        9'd484: Q <= 48'b000000000000000101110111000000000000101110001010;
        9'd485: Q <= 48'b000000000000100111110101000000000000001100001100;
        9'd486: Q <= 48'b000000000000100000101010000000000000010011010111;
        9'd487: Q <= 48'b000000000000011001101101000000000000011010010100;
        9'd488: Q <= 48'b000000000000010000100111000000000000100011011010;
        9'd489: Q <= 48'b000000000000000100111111000000000000101111000010;
        9'd490: Q <= 48'b000000000000101011010101000000000000001000101100;
        9'd491: Q <= 48'b000000000000001011110101000000000000101000001100;
        9'd492: Q <= 48'b000000000000100000110011000000000000010011001110;
        9'd493: Q <= 48'b000000000000001000110001000000000000101011010000;
        9'd494: Q <= 48'b000000000000100110100010000000000000001101011111;
        9'd495: Q <= 48'b000000000000101000100010000000000000001011011111;
        9'd496: Q <= 48'b000000000000101011110100000000000000001000001101;
        9'd497: Q <= 48'b000000000000010001000100000000000000100010111101;
        9'd498: Q <= 48'b000000000000000110010011000000000000101101101110;
        9'd499: Q <= 48'b000000000000010000000010000000000000100011111111;
        9'd500: Q <= 48'b000000000000010001110111000000000000100010001010;
        9'd501: Q <= 48'b000000000000100001100110000000000000010010011011;
        9'd502: Q <= 48'b000000000000101011010111000000000000001000101010;
        9'd503: Q <= 48'b000000000000001101110110000000000000100110001011;
        9'd504: Q <= 48'b000000000000011010111010000000000000011001000111;
        9'd505: Q <= 48'b000000000000010010111100000000000000100001000101;
        9'd506: Q <= 48'b000000000000011101010010000000000000010110101111;
        9'd507: Q <= 48'b000000000000010000000101000000000000100011111100;
        9'd508: Q <= 48'b000000000000100000111110000000000000010011000011;
        9'd509: Q <= 48'b000000000000101101110111000000000000000110001010;
        9'd510: Q <= 48'b000000000000001101110101000000000000100110001100;
        9'd511: Q <= 48'b000000000000100001101010000000000000010010010111;
        endcase end         
        end
`elsif OP2
    always@(posedge clk)
        begin
        if(REN == 1'b1) begin
        case(A)
        8'd0:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd1:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd2:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd3:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd4:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd5:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd6:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd7:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd8:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd9:   Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd10:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd11:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd12:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd13:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd14:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd15:  Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd16:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd17:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd18:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd19:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd20:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd21:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd22:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd23:  Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd24:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd25:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd26:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd27:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd28:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd29:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd30:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd31:  Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd32:  Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd33:  Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd34:  Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd35:  Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd36:  Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd37:  Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd38:  Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd39:  Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd40:  Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd41:  Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd42:  Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd43:  Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd44:  Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd45:  Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd46:  Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd47:  Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd48:  Q <= 96'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        8'd49:  Q <= 96'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        8'd50:  Q <= 96'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        8'd51:  Q <= 96'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        8'd52:  Q <= 96'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        8'd53:  Q <= 96'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        8'd54:  Q <= 96'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        8'd55:  Q <= 96'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        8'd56:  Q <= 96'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        8'd57:  Q <= 96'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        8'd58:  Q <= 96'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        8'd59:  Q <= 96'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        8'd60:  Q <= 96'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        8'd61:  Q <= 96'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        8'd62:  Q <= 96'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        8'd63:  Q <= 96'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        8'd64:  Q <= 96'b000100101000000100101000000100101000000100101000000100101000000100101000000100101000000100101000;
        8'd65:  Q <= 96'b100110001111100110001111100110001111100110001111100110001111100110001111100110001111100110001111;
        8'd66:  Q <= 96'b010100111011010100111011010100111011010100111011010100111011010100111011010100111011010100111011;
        8'd67:  Q <= 96'b010111000100010111000100010111000100010111000100010111000100010111000100010111000100010111000100;
        8'd68:  Q <= 96'b101111100110101111100110101111100110101111100110101111100110101111100110101111100110101111100110;
        8'd69:  Q <= 96'b000000111000000000111000000000111000000000111000000000111000000000111000000000111000000000111000;
        8'd70:  Q <= 96'b100011000000100011000000100011000000100011000000100011000000100011000000100011000000100011000000;
        8'd71:  Q <= 96'b010100110101010100110101010100110101010100110101010100110101010100110101010100110101010100110101;
        8'd72:  Q <= 96'b010110010010010110010010010110010010010110010010010110010010010110010010010110010010010110010010;
        8'd73:  Q <= 96'b100000101110100000101110100000101110100000101110100000101110100000101110100000101110100000101110;
        8'd74:  Q <= 96'b001000010111001000010111001000010111001000010111001000010111001000010111001000010111001000010111;
        8'd75:  Q <= 96'b101101000010101101000010101101000010101101000010101101000010101101000010101101000010101101000010;
        8'd76:  Q <= 96'b100101011001100101011001100101011001100101011001100101011001100101011001100101011001100101011001;
        8'd77:  Q <= 96'b101100111111101100111111101100111111101100111111101100111111101100111111101100111111101100111111;
        8'd78:  Q <= 96'b011110110110011110110110011110110110011110110110011110110110011110110110011110110110011110110110;
        8'd79:  Q <= 96'b001100110101001100110101001100110101001100110101001100110101001100110101001100110101001100110101;
        8'd80:  Q <= 96'b000100100001000100100001000100100001000100100001000101001011000101001011000101001011000101001011;
        8'd81:  Q <= 96'b110010110101110010110101110010110101110010110101011011011100011011011100011011011100011011011100;
        8'd82:  Q <= 96'b010010101101010010101101010010101101010010101101100100000000100100000000100100000000100100000000;
        8'd83:  Q <= 96'b100011100101100011100101100011100101100011100101100000000111100000000111100000000111100000000111;
        8'd84:  Q <= 96'b001010001010001010001010001010001010001010001010011110111001011110111001011110111001011110111001;
        8'd85:  Q <= 96'b100111010001100111010001100111010001100111010001001001111000001001111000001001111000001001111000;
        8'd86:  Q <= 96'b101100110001101100110001101100110001101100110001000000100001000000100001000000100001000000100001;
        8'd87:  Q <= 96'b010100101000010100101000010100101000010100101000011101111011011101111011011101111011011101111011;
        8'd88:  Q <= 96'b100100001111100100001111100100001111100100001111010110011011010110011011010110011011010110011011;
        8'd89:  Q <= 96'b001100100111001100100111001100100111001100100111000111000100000111000100000111000100000111000100;
        8'd90:  Q <= 96'b010110011110010110011110010110011110010110011110101100110100101100110100101100110100101100110100;
        8'd91:  Q <= 96'b010111111110010111111110010111111110010111111110100101100010100101100010100101100010100101100010;
        8'd92:  Q <= 96'b101001010111101001010111101001010111101001010111101000111001101000111001101000111001101000111001;
        8'd93:  Q <= 96'b010111001001010111001001010111001001010111001001001010001000001010001000001010001000001010001000;
        8'd94:  Q <= 96'b100110101010100110101010100110101010100110101010110000100110110000100110110000100110110000100110;
        8'd95:  Q <= 96'b010011001011010011001011010011001011010011001011001110001110001110001110001110001110001110001110;
        8'd96:  Q <= 96'b000000010001000000010001101011001001101011001001001001000111001001000111101001011001101001011001;
        8'd97:  Q <= 96'b011001100101011001100101001011010011001011010011100011110000100011110000010001001100010001001100;
        8'd98:  Q <= 96'b010110000001010110000001101001100110101001100110110011010001110011010001000011101001000011101001;
        8'd99:  Q <= 96'b001011110100001011110100100001101100100001101100101111000111101111000111101111101010101111101010;
        8'd100: Q <= 96'b011010100111011010100111011001110011011001110011101011100101101011100101011011111101011011111101;
        8'd101: Q <= 96'b011100110111011100110111001110111000001110111000010110110101010110110101101001111111101001111111;
        8'd102: Q <= 96'b001110101011001110101011100100000100100100000100100110000101100110000101100101010100100101010100;
        8'd103: Q <= 96'b001011011101001011011101100100100001100100100001000100001100000100001100001010000001001010000001;
        8'd104: Q <= 96'b011000110000011000110000100011111010100011111010011111110101011111110101110010010100110010010100;
        8'd105: Q <= 96'b000101110111000101110111100111110101100111110101100000101010100000101010011001101101011001101101;
        8'd106: Q <= 96'b010000100111010000100111000100111111000100111111101011010101101011010101001011110101001011110101;
        8'd107: Q <= 96'b100000110011100000110011001000110001001000110001100110100010100110100010101000100010101000100010;
        8'd108: Q <= 96'b101011110100101011110100010001000100010001000100000110010011000110010011010000000010010000000010;
        8'd109: Q <= 96'b010001110111010001110111100001100110100001100110101011010111101011010111001101110110001101110110;
        8'd110: Q <= 96'b011010111010011010111010010010111100010010111100011101010010011101010010010000000101010000000101;
        8'd111: Q <= 96'b100000111110100000111110101101110111101101110111001101110101001101110101100001101010100001101010;
        8'd112: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd113: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd114: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd115: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd116: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd117: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd118: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd119: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd120: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd121: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd122: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd123: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd124: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd125: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd126: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd127: Q <= 96'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        8'd128: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd129: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd130: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd131: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd132: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd133: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd134: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd135: Q <= 96'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        8'd136: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd137: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd138: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd139: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd140: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd141: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd142: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd143: Q <= 96'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        8'd144: Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd145: Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd146: Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd147: Q <= 96'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        8'd148: Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd149: Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd150: Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd151: Q <= 96'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        8'd152: Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd153: Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd154: Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd155: Q <= 96'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        8'd156: Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd157: Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd158: Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd159: Q <= 96'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        8'd160: Q <= 96'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        8'd161: Q <= 96'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        8'd162: Q <= 96'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        8'd163: Q <= 96'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        8'd164: Q <= 96'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        8'd165: Q <= 96'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        8'd166: Q <= 96'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        8'd167: Q <= 96'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        8'd168: Q <= 96'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        8'd169: Q <= 96'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        8'd170: Q <= 96'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        8'd171: Q <= 96'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        8'd172: Q <= 96'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        8'd173: Q <= 96'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        8'd174: Q <= 96'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        8'd175: Q <= 96'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        8'd176: Q <= 96'b001100110101001100110101001100110101001100110101001100110101001100110101001100110101001100110101;
        8'd177: Q <= 96'b011110110110011110110110011110110110011110110110011110110110011110110110011110110110011110110110;
        8'd178: Q <= 96'b101100111111101100111111101100111111101100111111101100111111101100111111101100111111101100111111;
        8'd179: Q <= 96'b100101011001100101011001100101011001100101011001100101011001100101011001100101011001100101011001;
        8'd180: Q <= 96'b101101000010101101000010101101000010101101000010101101000010101101000010101101000010101101000010;
        8'd181: Q <= 96'b001000010111001000010111001000010111001000010111001000010111001000010111001000010111001000010111;
        8'd182: Q <= 96'b100000101110100000101110100000101110100000101110100000101110100000101110100000101110100000101110;
        8'd183: Q <= 96'b010110010010010110010010010110010010010110010010010110010010010110010010010110010010010110010010;
        8'd184: Q <= 96'b010100110101010100110101010100110101010100110101010100110101010100110101010100110101010100110101;
        8'd185: Q <= 96'b100011000000100011000000100011000000100011000000100011000000100011000000100011000000100011000000;
        8'd186: Q <= 96'b000000111000000000111000000000111000000000111000000000111000000000111000000000111000000000111000;
        8'd187: Q <= 96'b101111100110101111100110101111100110101111100110101111100110101111100110101111100110101111100110;
        8'd188: Q <= 96'b010111000100010111000100010111000100010111000100010111000100010111000100010111000100010111000100;
        8'd189: Q <= 96'b010100111011010100111011010100111011010100111011010100111011010100111011010100111011010100111011;
        8'd190: Q <= 96'b100110001111100110001111100110001111100110001111100110001111100110001111100110001111100110001111;
        8'd191: Q <= 96'b000100101000000100101000000100101000000100101000000100101000000100101000000100101000000100101000;
        8'd192: Q <= 96'b001110001110001110001110001110001110001110001110010011001011010011001011010011001011010011001011;
        8'd193: Q <= 96'b110000100110110000100110110000100110110000100110100110101010100110101010100110101010100110101010;
        8'd194: Q <= 96'b001010001000001010001000001010001000001010001000010111001001010111001001010111001001010111001001;
        8'd195: Q <= 96'b101000111001101000111001101000111001101000111001101001010111101001010111101001010111101001010111;
        8'd196: Q <= 96'b100101100010100101100010100101100010100101100010010111111110010111111110010111111110010111111110;
        8'd197: Q <= 96'b101100110100101100110100101100110100101100110100010110011110010110011110010110011110010110011110;
        8'd198: Q <= 96'b000111000100000111000100000111000100000111000100001100100111001100100111001100100111001100100111;
        8'd199: Q <= 96'b010110011011010110011011010110011011010110011011100100001111100100001111100100001111100100001111;
        8'd200: Q <= 96'b011101111011011101111011011101111011011101111011010100101000010100101000010100101000010100101000;
        8'd201: Q <= 96'b000000100001000000100001000000100001000000100001101100110001101100110001101100110001101100110001;
        8'd202: Q <= 96'b001001111000001001111000001001111000001001111000100111010001100111010001100111010001100111010001;
        8'd203: Q <= 96'b011110111001011110111001011110111001011110111001001010001010001010001010001010001010001010001010;
        8'd204: Q <= 96'b100000000111100000000111100000000111100000000111100011100101100011100101100011100101100011100101;
        8'd205: Q <= 96'b100100000000100100000000100100000000100100000000010010101101010010101101010010101101010010101101;
        8'd206: Q <= 96'b011011011100011011011100011011011100011011011100110010110101110010110101110010110101110010110101;
        8'd207: Q <= 96'b000101001011000101001011000101001011000101001011000100100001000100100001000100100001000100100001;
        8'd208: Q <= 96'b100001101010100001101010001101110101001101110101101101110111101101110111100000111110100000111110;
        8'd209: Q <= 96'b010000000101010000000101011101010010011101010010010010111100010010111100011010111010011010111010;
        8'd210: Q <= 96'b001101110110001101110110101011010111101011010111100001100110100001100110010001110111010001110111;
        8'd211: Q <= 96'b010000000010010000000010000110010011000110010011010001000100010001000100101011110100101011110100;
        8'd212: Q <= 96'b101000100010101000100010100110100010100110100010001000110001001000110001100000110011100000110011;
        8'd213: Q <= 96'b001011110101001011110101101011010101101011010101000100111111000100111111010000100111010000100111;
        8'd214: Q <= 96'b011001101101011001101101100000101010100000101010100111110101100111110101000101110111000101110111;
        8'd215: Q <= 96'b110010010100110010010100011111110101011111110101100011111010100011111010011000110000011000110000;
        8'd216: Q <= 96'b001010000001001010000001000100001100000100001100100100100001100100100001001011011101001011011101;
        8'd217: Q <= 96'b100101010100100101010100100110000101100110000101100100000100100100000100001110101011001110101011;
        8'd218: Q <= 96'b101001111111101001111111010110110101010110110101001110111000001110111000011100110111011100110111;
        8'd219: Q <= 96'b011011111101011011111101101011100101101011100101011001110011011001110011011010100111011010100111;
        8'd220: Q <= 96'b101111101010101111101010101111000111101111000111100001101100100001101100001011110100001011110100;
        8'd221: Q <= 96'b000011101001000011101001110011010001110011010001101001100110101001100110010110000001010110000001;
        8'd222: Q <= 96'b010001001100010001001100100011110000100011110000001011010011001011010011011001100101011001100101;
        8'd223: Q <= 96'b101001011001101001011001001001000111001001000111101011001001101011001001000000010001000000010001;
        8'd224: Q <= 96'b000000000000000000010001000000000000110011110000000000000000101011001001000000000000001000111000;
        8'd225: Q <= 96'b000000000000001001000111000000000000101010111010000000000000101001011001000000000000001010101000;
        8'd226: Q <= 96'b000000000000011001100101000000000000011010011100000000000000001011010011000000000000101000101110;
        8'd227: Q <= 96'b000000000000100011110000000000000000010000010001000000000000010001001100000000000000100010110101;
        8'd228: Q <= 96'b000000000000010110000001000000000000011110000000000000000000101001100110000000000000001010011011;
        8'd229: Q <= 96'b000000000000110011010001000000000000000000110000000000000000000011101001000000000000110000011000;
        8'd230: Q <= 96'b000000000000001011110100000000000000101000001101000000000000100001101100000000000000010010010101;
        8'd231: Q <= 96'b000000000000101111000111000000000000000100111010000000000000101111101010000000000000000100010111;
        8'd232: Q <= 96'b000000000000011010100111000000000000011001011010000000000000011001110011000000000000011010001110;
        8'd233: Q <= 96'b000000000000101011100101000000000000001000011100000000000000011011111101000000000000011000000100;
        8'd234: Q <= 96'b000000000000011100110111000000000000010111001010000000000000001110111000000000000000100101001001;
        8'd235: Q <= 96'b000000000000010110110101000000000000011101001100000000000000101001111111000000000000001010000010;
        8'd236: Q <= 96'b000000000000001110101011000000000000100101010110000000000000100100000100000000000000001111111101;
        8'd237: Q <= 96'b000000000000100110000101000000000000001101111100000000000000100101010100000000000000001110101101;
        8'd238: Q <= 96'b000000000000001011011101000000000000101000100100000000000000100100100001000000000000001111100000;
        8'd239: Q <= 96'b000000000000000100001100000000000000101111110101000000000000001010000001000000000000101010000000;
        8'd240: Q <= 96'b000000000000011000110000000000000000011011010001000000000000100011111010000000000000010000000111;
        8'd241: Q <= 96'b000000000000011111110101000000000000010100001100000000000000110010010100000000000000000001101101;
        8'd242: Q <= 96'b000000000000000101110111000000000000101110001010000000000000100111110101000000000000001100001100;
        8'd243: Q <= 96'b000000000000100000101010000000000000010011010111000000000000011001101101000000000000011010010100;
        8'd244: Q <= 96'b000000000000010000100111000000000000100011011010000000000000000100111111000000000000101111000010;
        8'd245: Q <= 96'b000000000000101011010101000000000000001000101100000000000000001011110101000000000000101000001100;
        8'd246: Q <= 96'b000000000000100000110011000000000000010011001110000000000000001000110001000000000000101011010000;
        8'd247: Q <= 96'b000000000000100110100010000000000000001101011111000000000000101000100010000000000000001011011111;
        8'd248: Q <= 96'b000000000000101011110100000000000000001000001101000000000000010001000100000000000000100010111101;
        8'd249: Q <= 96'b000000000000000110010011000000000000101101101110000000000000010000000010000000000000100011111111;
        8'd250: Q <= 96'b000000000000010001110111000000000000100010001010000000000000100001100110000000000000010010011011;
        8'd251: Q <= 96'b000000000000101011010111000000000000001000101010000000000000001101110110000000000000100110001011;
        8'd252: Q <= 96'b000000000000011010111010000000000000011001000111000000000000010010111100000000000000100001000101;
        8'd253: Q <= 96'b000000000000011101010010000000000000010110101111000000000000010000000101000000000000100011111100;
        8'd254: Q <= 96'b000000000000100000111110000000000000010011000011000000000000101101110111000000000000000110001010;
        8'd255: Q <= 96'b000000000000001101110101000000000000100110001100000000000000100001101010000000000000010010010111;
        endcase end         
        end
`else 
    always@(posedge clk)
        begin
        if(REN == 1'b1) begin
        case(A)
        7'd0:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd1:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd2:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd3:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd4:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd5:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd6:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd7:   Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd8:   Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd9:   Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd10:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd11:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd12:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd13:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd14:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd15:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd16:  Q<=192'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        7'd17:  Q<=192'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        7'd18:  Q<=192'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        7'd19:  Q<=192'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        7'd20:  Q<=192'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        7'd21:  Q<=192'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        7'd22:  Q<=192'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        7'd23:  Q<=192'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        7'd24:  Q<=192'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        7'd25:  Q<=192'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        7'd26:  Q<=192'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        7'd27:  Q<=192'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        7'd28:  Q<=192'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        7'd29:  Q<=192'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        7'd30:  Q<=192'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        7'd31:  Q<=192'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        7'd32:  Q<=192'b000100101000000100101000000100101000000100101000000100101000000100101000000100101000000100101000100110001111100110001111100110001111100110001111100110001111100110001111100110001111100110001111;
        7'd33:  Q<=192'b010100111011010100111011010100111011010100111011010100111011010100111011010100111011010100111011010111000100010111000100010111000100010111000100010111000100010111000100010111000100010111000100;
        7'd34:  Q<=192'b101111100110101111100110101111100110101111100110101111100110101111100110101111100110101111100110000000111000000000111000000000111000000000111000000000111000000000111000000000111000000000111000;
        7'd35:  Q<=192'b100011000000100011000000100011000000100011000000100011000000100011000000100011000000100011000000010100110101010100110101010100110101010100110101010100110101010100110101010100110101010100110101;
        7'd36:  Q<=192'b010110010010010110010010010110010010010110010010010110010010010110010010010110010010010110010010100000101110100000101110100000101110100000101110100000101110100000101110100000101110100000101110;
        7'd37:  Q<=192'b001000010111001000010111001000010111001000010111001000010111001000010111001000010111001000010111101101000010101101000010101101000010101101000010101101000010101101000010101101000010101101000010;
        7'd38:  Q<=192'b100101011001100101011001100101011001100101011001100101011001100101011001100101011001100101011001101100111111101100111111101100111111101100111111101100111111101100111111101100111111101100111111;
        7'd39:  Q<=192'b011110110110011110110110011110110110011110110110011110110110011110110110011110110110011110110110001100110101001100110101001100110101001100110101001100110101001100110101001100110101001100110101;
        7'd40:  Q<=192'b000100100001000100100001000100100001000100100001000101001011000101001011000101001011000101001011110010110101110010110101110010110101110010110101011011011100011011011100011011011100011011011100;
        7'd41:  Q<=192'b010010101101010010101101010010101101010010101101100100000000100100000000100100000000100100000000100011100101100011100101100011100101100011100101100000000111100000000111100000000111100000000111;
        7'd42:  Q<=192'b001010001010001010001010001010001010001010001010011110111001011110111001011110111001011110111001100111010001100111010001100111010001100111010001001001111000001001111000001001111000001001111000;
        7'd43:  Q<=192'b101100110001101100110001101100110001101100110001000000100001000000100001000000100001000000100001010100101000010100101000010100101000010100101000011101111011011101111011011101111011011101111011;
        7'd44:  Q<=192'b100100001111100100001111100100001111100100001111010110011011010110011011010110011011010110011011001100100111001100100111001100100111001100100111000111000100000111000100000111000100000111000100;
        7'd45:  Q<=192'b010110011110010110011110010110011110010110011110101100110100101100110100101100110100101100110100010111111110010111111110010111111110010111111110100101100010100101100010100101100010100101100010;
        7'd46:  Q<=192'b101001010111101001010111101001010111101001010111101000111001101000111001101000111001101000111001010111001001010111001001010111001001010111001001001010001000001010001000001010001000001010001000;
        7'd47:  Q<=192'b100110101010100110101010100110101010100110101010110000100110110000100110110000100110110000100110010011001011010011001011010011001011010011001011001110001110001110001110001110001110001110001110;
        7'd48:  Q<=192'b000000010001000000010001101011001001101011001001001001000111001001000111101001011001101001011001011001100101011001100101001011010011001011010011100011110000100011110000010001001100010001001100;
        7'd49:  Q<=192'b010110000001010110000001101001100110101001100110110011010001110011010001000011101001000011101001001011110100001011110100100001101100100001101100101111000111101111000111101111101010101111101010;
        7'd50:  Q<=192'b011010100111011010100111011001110011011001110011101011100101101011100101011011111101011011111101011100110111011100110111001110111000001110111000010110110101010110110101101001111111101001111111;
        7'd51:  Q<=192'b001110101011001110101011100100000100100100000100100110000101100110000101100101010100100101010100001011011101001011011101100100100001100100100001000100001100000100001100001010000001001010000001;
        7'd52:  Q<=192'b011000110000011000110000100011111010100011111010011111110101011111110101110010010100110010010100000101110111000101110111100111110101100111110101100000101010100000101010011001101101011001101101;
        7'd53:  Q<=192'b010000100111010000100111000100111111000100111111101011010101101011010101001011110101001011110101100000110011100000110011001000110001001000110001100110100010100110100010101000100010101000100010;
        7'd54:  Q<=192'b101011110100101011110100010001000100010001000100000110010011000110010011010000000010010000000010010001110111010001110111100001100110100001100110101011010111101011010111001101110110001101110110;
        7'd55:  Q<=192'b011010111010011010111010010010111100010010111100011101010010011101010010010000000101010000000101100000111110100000111110101101110111101101110111001101110101001101110101100001101010100001101010;
        7'd56:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd57:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd58:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd59:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd60:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd61:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd62:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd63:  Q<=192'b011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001011011000001;
        7'd64:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd65:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd66:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd67:  Q<=192'b110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001110011011001;
        7'd68:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd69:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd70:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd71:  Q<=192'b101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100101000010100;
        7'd72:  Q<=192'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        7'd73:  Q<=192'b001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000001101010000;
        7'd74:  Q<=192'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        7'd75:  Q<=192'b011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001011101101001;
        7'd76:  Q<=192'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        7'd77:  Q<=192'b001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110001001110110;
        7'd78:  Q<=192'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        7'd79:  Q<=192'b101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010101001010010;
        7'd80:  Q<=192'b011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010011011010010;
        7'd81:  Q<=192'b001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001001000111001;
        7'd82:  Q<=192'b110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100110010111100;
        7'd83:  Q<=192'b101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010101011100010;
        7'd84:  Q<=192'b001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101001100011101;
        7'd85:  Q<=192'b000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001000011000001;
        7'd86:  Q<=192'b011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111011101111111;
        7'd87:  Q<=192'b010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110010000100110;
        7'd88:  Q<=192'b001100110101001100110101001100110101001100110101001100110101001100110101001100110101001100110101011110110110011110110110011110110110011110110110011110110110011110110110011110110110011110110110;
        7'd89:  Q<=192'b101100111111101100111111101100111111101100111111101100111111101100111111101100111111101100111111100101011001100101011001100101011001100101011001100101011001100101011001100101011001100101011001;
        7'd90:  Q<=192'b101101000010101101000010101101000010101101000010101101000010101101000010101101000010101101000010001000010111001000010111001000010111001000010111001000010111001000010111001000010111001000010111;
        7'd91:  Q<=192'b100000101110100000101110100000101110100000101110100000101110100000101110100000101110100000101110010110010010010110010010010110010010010110010010010110010010010110010010010110010010010110010010;
        7'd92:  Q<=192'b010100110101010100110101010100110101010100110101010100110101010100110101010100110101010100110101100011000000100011000000100011000000100011000000100011000000100011000000100011000000100011000000;
        7'd93:  Q<=192'b000000111000000000111000000000111000000000111000000000111000000000111000000000111000000000111000101111100110101111100110101111100110101111100110101111100110101111100110101111100110101111100110;
        7'd94:  Q<=192'b010111000100010111000100010111000100010111000100010111000100010111000100010111000100010111000100010100111011010100111011010100111011010100111011010100111011010100111011010100111011010100111011;
        7'd95:  Q<=192'b100110001111100110001111100110001111100110001111100110001111100110001111100110001111100110001111000100101000000100101000000100101000000100101000000100101000000100101000000100101000000100101000;
        7'd96:  Q<=192'b001110001110001110001110001110001110001110001110010011001011010011001011010011001011010011001011110000100110110000100110110000100110110000100110100110101010100110101010100110101010100110101010;
        7'd97:  Q<=192'b001010001000001010001000001010001000001010001000010111001001010111001001010111001001010111001001101000111001101000111001101000111001101000111001101001010111101001010111101001010111101001010111;
        7'd98:  Q<=192'b100101100010100101100010100101100010100101100010010111111110010111111110010111111110010111111110101100110100101100110100101100110100101100110100010110011110010110011110010110011110010110011110;
        7'd99:  Q<=192'b000111000100000111000100000111000100000111000100001100100111001100100111001100100111001100100111010110011011010110011011010110011011010110011011100100001111100100001111100100001111100100001111;
        7'd100: Q<=192'b011101111011011101111011011101111011011101111011010100101000010100101000010100101000010100101000000000100001000000100001000000100001000000100001101100110001101100110001101100110001101100110001;
        7'd101: Q<=192'b001001111000001001111000001001111000001001111000100111010001100111010001100111010001100111010001011110111001011110111001011110111001011110111001001010001010001010001010001010001010001010001010;
        7'd102: Q<=192'b100000000111100000000111100000000111100000000111100011100101100011100101100011100101100011100101100100000000100100000000100100000000100100000000010010101101010010101101010010101101010010101101;
        7'd103: Q<=192'b011011011100011011011100011011011100011011011100110010110101110010110101110010110101110010110101000101001011000101001011000101001011000101001011000100100001000100100001000100100001000100100001;
        7'd104: Q<=192'b100001101010100001101010001101110101001101110101101101110111101101110111100000111110100000111110010000000101010000000101011101010010011101010010010010111100010010111100011010111010011010111010;
        7'd105: Q<=192'b001101110110001101110110101011010111101011010111100001100110100001100110010001110111010001110111010000000010010000000010000110010011000110010011010001000100010001000100101011110100101011110100;
        7'd106: Q<=192'b101000100010101000100010100110100010100110100010001000110001001000110001100000110011100000110011001011110101001011110101101011010101101011010101000100111111000100111111010000100111010000100111;
        7'd107: Q<=192'b011001101101011001101101100000101010100000101010100111110101100111110101000101110111000101110111110010010100110010010100011111110101011111110101100011111010100011111010011000110000011000110000;
        7'd108: Q<=192'b001010000001001010000001000100001100000100001100100100100001100100100001001011011101001011011101100101010100100101010100100110000101100110000101100100000100100100000100001110101011001110101011;
        7'd109: Q<=192'b101001111111101001111111010110110101010110110101001110111000001110111000011100110111011100110111011011111101011011111101101011100101101011100101011001110011011001110011011010100111011010100111;
        7'd110: Q<=192'b101111101010101111101010101111000111101111000111100001101100100001101100001011110100001011110100000011101001000011101001110011010001110011010001101001100110101001100110010110000001010110000001;
        7'd111: Q<=192'b010001001100010001001100100011110000100011110000001011010011001011010011011001100101011001100101101001011001101001011001001001000111001001000111101011001001101011001001000000010001000000010001;
        7'd112: Q<=192'b000000000000000000010001000000000000110011110000000000000000101011001001000000000000001000111000000000000000001001000111000000000000101010111010000000000000101001011001000000000000001010101000;
        7'd113: Q<=192'b000000000000011001100101000000000000011010011100000000000000001011010011000000000000101000101110000000000000100011110000000000000000010000010001000000000000010001001100000000000000100010110101;
        7'd114: Q<=192'b000000000000010110000001000000000000011110000000000000000000101001100110000000000000001010011011000000000000110011010001000000000000000000110000000000000000000011101001000000000000110000011000;
        7'd115: Q<=192'b000000000000001011110100000000000000101000001101000000000000100001101100000000000000010010010101000000000000101111000111000000000000000100111010000000000000101111101010000000000000000100010111;
        7'd116: Q<=192'b000000000000011010100111000000000000011001011010000000000000011001110011000000000000011010001110000000000000101011100101000000000000001000011100000000000000011011111101000000000000011000000100;
        7'd117: Q<=192'b000000000000011100110111000000000000010111001010000000000000001110111000000000000000100101001001000000000000010110110101000000000000011101001100000000000000101001111111000000000000001010000010;
        7'd118: Q<=192'b000000000000001110101011000000000000100101010110000000000000100100000100000000000000001111111101000000000000100110000101000000000000001101111100000000000000100101010100000000000000001110101101;
        7'd119: Q<=192'b000000000000001011011101000000000000101000100100000000000000100100100001000000000000001111100000000000000000000100001100000000000000101111110101000000000000001010000001000000000000101010000000;
        7'd120: Q<=192'b000000000000011000110000000000000000011011010001000000000000100011111010000000000000010000000111000000000000011111110101000000000000010100001100000000000000110010010100000000000000000001101101;
        7'd121: Q<=192'b000000000000000101110111000000000000101110001010000000000000100111110101000000000000001100001100000000000000100000101010000000000000010011010111000000000000011001101101000000000000011010010100;
        7'd122: Q<=192'b000000000000010000100111000000000000100011011010000000000000000100111111000000000000101111000010000000000000101011010101000000000000001000101100000000000000001011110101000000000000101000001100;
        7'd123: Q<=192'b000000000000100000110011000000000000010011001110000000000000001000110001000000000000101011010000000000000000100110100010000000000000001101011111000000000000101000100010000000000000001011011111;
        7'd124: Q<=192'b000000000000101011110100000000000000001000001101000000000000010001000100000000000000100010111101000000000000000110010011000000000000101101101110000000000000010000000010000000000000100011111111;
        7'd125: Q<=192'b000000000000010001110111000000000000100010001010000000000000100001100110000000000000010010011011000000000000101011010111000000000000001000101010000000000000001101110110000000000000100110001011;
        7'd126: Q<=192'b000000000000011010111010000000000000011001000111000000000000010010111100000000000000100001000101000000000000011101010010000000000000010110101111000000000000010000000101000000000000100011111100;
        7'd127: Q<=192'b000000000000100000111110000000000000010011000011000000000000101101110111000000000000000110001010000000000000001101110101000000000000100110001100000000000000100001101010000000000000010010010111;
        endcase end         
        end
`endif

endmodule