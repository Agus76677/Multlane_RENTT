`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: HZW
// 
// Create Date: 2025/03/28 18:32:12
// Design Name: 
// Module Name: Hybrid_compress_Red_wocsa3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// Modulus by bit
module Hybrid_compress_Red_wocsa3(
    input [8-1:0] t0_0,
    input [4-1:0] t0_1,
    input [6-1:0] t0_2,
    input [5-1:0] t0_3,
    input [4-1:0] t0_4,
    input [5-1:0] t0_5,
    input [5-1:0] t0_6,
    input [4-1:0] t0_7,
    input [5-1:0] t0_8,
    input [6-1:0] t0_9,
    input [6-1:0] t0_10,
    input [1-1:0] t0_11,
    // input [1-1:0] t0_12,
    // input [1-1:0] t0_13,
    // input [1-1:0] t0_14,
    output [14-1:0] s,
    output [15-1:0] c);

// ------------------------------- Connections
    // --------------------- Level 1
    wire [4-1:0] t1_0;
    wire [4-1:0] t1_1;
    wire [4-1:0] t1_2;
    wire [4-1:0] t1_3;
    wire [4-1:0] t1_4;
    wire [4-1:0] t1_5;
    wire [4-1:0] t1_6;
    wire [4-1:0] t1_7;
    wire [4-1:0] t1_8;
    wire [4-1:0] t1_9;
    wire [4-1:0] t1_10;
    wire [3-1:0] t1_11;
    // wire [1-1:0] t1_12;
    // wire [1-1:0] t1_13;
    // wire [1-1:0] t1_14;

    // --------------------- Level 2
    wire [2-1:0] t2_0;
    wire [3-1:0] t2_1;
    wire [3-1:0] t2_2;
    wire [3-1:0] t2_3;
    wire [3-1:0] t2_4;
    wire [3-1:0] t2_5;
    wire [3-1:0] t2_6;
    wire [3-1:0] t2_7;
    wire [3-1:0] t2_8;
    wire [3-1:0] t2_9;
    wire [3-1:0] t2_10;
    wire [2-1:0] t2_11;
    wire [1-1:0] t2_12;
    // wire [2-1:0] t2_12;
    // wire [1-1:0] t2_13;
    // wire [1-1:0] t2_14;

    // --------------------- Level 3
    wire [2-1:0] t3_0;
    wire [2-1:0] t3_1;
    wire [2-1:0] t3_2;
    wire [2-1:0] t3_3;
    wire [2-1:0] t3_4;
    wire [2-1:0] t3_5;
    wire [2-1:0] t3_6;
    wire [2-1:0] t3_7;
    wire [2-1:0] t3_8;
    wire [2-1:0] t3_9;
    wire [2-1:0] t3_10;
    wire [2-1:0] t3_11;
    wire [2-1:0] t3_12;
    wire [1-1:0] t3_13;
    // wire [2-1:0] t3_13;
    // wire [1-1:0] t3_14;
// ------------------------------- Operations

    // --------------------- Level 1
    // 0
    // CSA3 u000(t0_0[0],t0_0[1],t0_0[2],t0_0[3],t0_0[4],t1_0[0],t1_1[0],t1_1[1]);
    CSA2 u000(t0_0[0],t0_0[1],t0_0[2],t1_0[0],t1_1[0]);
    CSA2 u001(t0_0[3],t0_0[4],t0_0[5],t1_0[1],t1_1[1]);
    // assign t1_0[1] = t0_0[5];
    assign t1_0[2] = t0_0[6];
    assign t1_0[3] = t0_0[7];
    // 1
    CSA2 u010(t0_1[0],t0_1[1],t0_1[2],t1_1[2],t1_2[0]);
    assign t1_1[3] = t0_1[3];
    // 2
    CSA2 u020(t0_2[0],t0_2[1],t0_2[2],t1_2[1],t1_3[0]);
    CSA1 u021(t0_2[3],t0_2[4],t1_2[2],t1_3[1]);
    assign t1_2[3] = t0_2[5];
    // 3
    CSA2 u030(t0_3[0],t0_3[1],t0_3[2],t1_3[2],t1_4[0]);
    CSA1 u031(t0_3[3],t0_3[4],t1_3[3],t1_4[1]);
    // 4
    CSA2 u040(t0_4[0],t0_4[1],t0_4[2],t1_4[2],t1_5[0]);
    assign t1_4[3] = t0_4[3];
    // 5
    CSA2 u050(t0_5[0],t0_5[1],t0_5[2],t1_5[1],t1_6[0]);
    assign t1_5[2] = t0_5[3];
    assign t1_5[3] = t0_5[4];
    // 6
    CSA2 u060(t0_6[0],t0_6[1],t0_6[2],t1_6[1],t1_7[0]);
    assign t1_6[2] = t0_6[3];
    assign t1_6[3] = t0_6[4];
  
    // 7
    CSA1 u070(t0_7[0],t0_7[1],t1_7[1],t1_8[0]);
    assign t1_7[2] = t0_7[2];
    assign t1_7[3] = t0_7[3];
    // 8
    CSA2 u080(t0_8[0],t0_8[1],t0_8[2],t1_8[1],t1_9[0]);
    assign t1_8[2] = t0_8[3];
    assign t1_8[3] = t0_8[4];
    
    // 9
    CSA2 u090(t0_9[0],t0_9[1],t0_9[2],t1_9[1],t1_10[0]);
    CSA1 u091(t0_9[3],t0_9[4],t1_9[2],t1_10[1]);
    assign t1_9[3] = t0_9[5];

    // 10
    CSA2 u0100(t0_10[0],t0_10[1],t0_10[2],t1_10[2],t1_11[0]);
    CSA2 u0101(t0_10[3],t0_10[4],t0_10[5],t1_10[3],t1_11[1]);

    assign t1_11[2] = t0_11[0];
    // assign t1_12[0] = t0_12[0];
    // assign t1_13[0] = t0_13[0];
    // assign t1_14[0] = t0_14[0];

    // --------------------- Level 2
    // 0
    CSA2 u100(t1_0[0],t1_0[1],t1_0[2],t2_0[0],t2_1[0]);
    assign t2_0[1] = t1_0[3];
    // 1
    CSA2 u110(t1_1[0],t1_1[1],t1_1[2],t2_1[1],t2_2[0]);
    assign t2_1[2] = t1_1[3];
    // 2
    CSA2 u120(t1_2[0],t1_2[1],t1_2[2],t2_2[1],t2_3[0]);
    assign t2_2[2] = t1_2[3];
    // 3
    CSA2 u130(t1_3[0],t1_3[1],t1_3[2],t2_3[1],t2_4[0]);
    assign t2_3[2] = t1_3[3];
    // 4   
    CSA2 u140(t1_4[0],t1_4[1],t1_4[2],t2_4[1],t2_5[0]);
    assign t2_4[2] = t1_4[3];
    // 5
    CSA2 u150(t1_5[0],t1_5[1],t1_5[2],t2_5[1],t2_6[0]);
    assign t2_5[2] = t1_5[3];
    // 6
    CSA2 u160(t1_6[0],t1_6[1],t1_6[2],t2_6[1],t2_7[0]);
    assign t2_6[2] = t1_6[3];
    // 7
    CSA2 u170(t1_7[0],t1_7[1],t1_7[2],t2_7[1],t2_8[0]);
    assign t2_7[2] = t1_7[3];
    // 8    
    CSA2 u180(t1_8[0],t1_8[1],t1_8[2],t2_8[1],t2_9[0]);
    assign t2_8[2] = t1_8[3];
    // 9
    CSA2 u190(t1_9[0],t1_9[1],t1_9[2],t2_9[1],t2_10[0]); 
    assign t2_9[2] = t1_9[3];
    // 10
    CSA2 u1100(t1_10[0],t1_10[1],t1_10[2],t2_10[1],t2_11[0]);
    assign t2_10[2] = t1_10[3];
    // 11
    CSA2 u1110(t1_11[0],t1_11[1],t1_11[2],t2_11[1],t2_12[0]);
    // assign t2_12[1] = 1'b1;

    // assign t2_12[1] = t1_12[0];
    // assign t2_13[0] = t1_13[0];
    // assign t2_14[0] = t1_14[0];

    // --------------------- Level 3
    // 0
    assign t3_0[0] = t2_0[0];
    assign t3_0[1] = t2_0[1];
    // 1
    CSA1 u21(t2_1[0],t2_1[1],t3_1[0],t3_2[0]);
    assign t3_1[1] = t2_1[2];
    // 2
    CSA2 u22(t2_2[0],t2_2[1],t2_2[2],t3_2[1],t3_3[0]);
    // 3
    CSA2 u23(t2_3[0],t2_3[1],t2_3[2],t3_3[1],t3_4[0]);
    // 4
    CSA2 u24(t2_4[0],t2_4[1],t2_4[2],t3_4[1],t3_5[0]);
    // 5
    CSA2 u25(t2_5[0],t2_5[1],t2_5[2],t3_5[1],t3_6[0]);
    // 6
    CSA2 u26(t2_6[0],t2_6[1],t2_6[2],t3_6[1],t3_7[0]);
    // 7 
    CSA2 u27(t2_7[0],t2_7[1],t2_7[2],t3_7[1],t3_8[0]);
    // 8
    CSA2 u28(t2_8[0],t2_8[1],t2_8[2],t3_8[1],t3_9[0]);
    // 9
    CSA2 u29(t2_9[0],t2_9[1],t2_9[2],t3_9[1],t3_10[0]);
    // 10
    CSA2 u210(t2_10[0],t2_10[1],t2_10[2],t3_10[1],t3_11[0]);
    // 11
    CSA1 u211(t2_11[0],t2_11[1],t3_11[1],t3_12[0]);
    // 12
    CSA1 u212(t2_12[0],1'b1,t3_12[1],t3_13[0]);

    // assign t3_13[1] = 1'b1;
    // assign t3_14[0] = 1'b1;


    // assign t3_13[1] = t2_13[0];
    // assign t3_14[0] = t2_14[0];

    // --------------------- Rewire

    assign c[0]  = t3_0[0];
    assign c[1]  = t3_1[0];
    assign c[2]  = t3_2[0];
    assign c[3]  = t3_3[0];
    assign c[4]  = t3_4[0];
    assign c[5]  = t3_5[0];
    assign c[6]  = t3_6[0];
    assign c[7]  = t3_7[0];
    assign c[8]  = t3_8[0];
    assign c[9]  = t3_9[0];
    assign c[10] = t3_10[0];
    assign c[11] = t3_11[0];
    assign c[12] = t3_12[0];
    assign c[13] = t3_13[0];
    assign c[14] = 1'b1;
    assign s[0]  = t3_0[1];
    assign s[1]  = t3_1[1];
    assign s[2]  = t3_2[1];
    assign s[3]  = t3_3[1];
    assign s[4]  = t3_4[1];
    assign s[5]  = t3_5[1];
    assign s[6]  = t3_6[1];
    assign s[7]  = t3_7[1];
    assign s[8]  = t3_8[1];
    assign s[9]  = t3_9[1];
    assign s[10] = t3_10[1];
    assign s[11] = t3_11[1];
    assign s[12] = t3_12[1];
    assign s[13] = 1'b1;
    // assign s[14] = 1'b0;

endmodule